// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 15.0.0 Build 145 04/22/2015 SJ Full Version"

// DATE "07/12/2016 09:11:56"

// 
// Device: Altera 5CSEMA5F31C6 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module NCO_Lab3 (
	clk,
	clken,
	phi_inc_i,
	fsin_o,
	out_valid,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	clken;
input 	[31:0] phi_inc_i;
output 	[11:0] fsin_o;
output 	out_valid;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nco_ii_0|sop|sin_o[0]~q ;
wire \nco_ii_0|sop|sin_o[1]~q ;
wire \nco_ii_0|sop|sin_o[2]~q ;
wire \nco_ii_0|sop|sin_o[3]~q ;
wire \nco_ii_0|sop|sin_o[4]~q ;
wire \nco_ii_0|sop|sin_o[5]~q ;
wire \nco_ii_0|sop|sin_o[6]~q ;
wire \nco_ii_0|sop|sin_o[7]~q ;
wire \nco_ii_0|sop|sin_o[8]~q ;
wire \nco_ii_0|sop|sin_o[9]~q ;
wire \nco_ii_0|sop|sin_o[10]~q ;
wire \nco_ii_0|sop|sin_o[11]~q ;
wire \nco_ii_0|ux710isdr|data_ready~q ;
wire \clk~input_o ;
wire \reset_n~input_o ;
wire \clken~input_o ;
wire \phi_inc_i[30]~input_o ;
wire \phi_inc_i[31]~input_o ;
wire \phi_inc_i[29]~input_o ;
wire \phi_inc_i[28]~input_o ;
wire \phi_inc_i[27]~input_o ;
wire \phi_inc_i[26]~input_o ;
wire \phi_inc_i[25]~input_o ;
wire \phi_inc_i[24]~input_o ;
wire \phi_inc_i[23]~input_o ;
wire \phi_inc_i[22]~input_o ;
wire \phi_inc_i[21]~input_o ;
wire \phi_inc_i[20]~input_o ;
wire \phi_inc_i[19]~input_o ;
wire \phi_inc_i[18]~input_o ;
wire \phi_inc_i[17]~input_o ;
wire \phi_inc_i[16]~input_o ;
wire \phi_inc_i[15]~input_o ;
wire \phi_inc_i[14]~input_o ;
wire \phi_inc_i[13]~input_o ;
wire \phi_inc_i[12]~input_o ;
wire \phi_inc_i[11]~input_o ;
wire \phi_inc_i[10]~input_o ;
wire \phi_inc_i[9]~input_o ;
wire \phi_inc_i[8]~input_o ;
wire \phi_inc_i[7]~input_o ;
wire \phi_inc_i[6]~input_o ;
wire \phi_inc_i[5]~input_o ;
wire \phi_inc_i[4]~input_o ;
wire \phi_inc_i[3]~input_o ;
wire \phi_inc_i[2]~input_o ;
wire \phi_inc_i[1]~input_o ;
wire \phi_inc_i[0]~input_o ;


NCO_Lab3_NCO_Lab3_nco_ii_0 nco_ii_0(
	.sin_o_0(\nco_ii_0|sop|sin_o[0]~q ),
	.sin_o_1(\nco_ii_0|sop|sin_o[1]~q ),
	.sin_o_2(\nco_ii_0|sop|sin_o[2]~q ),
	.sin_o_3(\nco_ii_0|sop|sin_o[3]~q ),
	.sin_o_4(\nco_ii_0|sop|sin_o[4]~q ),
	.sin_o_5(\nco_ii_0|sop|sin_o[5]~q ),
	.sin_o_6(\nco_ii_0|sop|sin_o[6]~q ),
	.sin_o_7(\nco_ii_0|sop|sin_o[7]~q ),
	.sin_o_8(\nco_ii_0|sop|sin_o[8]~q ),
	.sin_o_9(\nco_ii_0|sop|sin_o[9]~q ),
	.sin_o_10(\nco_ii_0|sop|sin_o[10]~q ),
	.sin_o_11(\nco_ii_0|sop|sin_o[11]~q ),
	.data_ready(\nco_ii_0|ux710isdr|data_ready~q ),
	.clk(\clk~input_o ),
	.reset_n(\reset_n~input_o ),
	.clken(\clken~input_o ),
	.phi_inc_i_30(\phi_inc_i[30]~input_o ),
	.phi_inc_i_31(\phi_inc_i[31]~input_o ),
	.phi_inc_i_29(\phi_inc_i[29]~input_o ),
	.phi_inc_i_28(\phi_inc_i[28]~input_o ),
	.phi_inc_i_27(\phi_inc_i[27]~input_o ),
	.phi_inc_i_26(\phi_inc_i[26]~input_o ),
	.phi_inc_i_25(\phi_inc_i[25]~input_o ),
	.phi_inc_i_24(\phi_inc_i[24]~input_o ),
	.phi_inc_i_23(\phi_inc_i[23]~input_o ),
	.phi_inc_i_22(\phi_inc_i[22]~input_o ),
	.phi_inc_i_21(\phi_inc_i[21]~input_o ),
	.phi_inc_i_20(\phi_inc_i[20]~input_o ),
	.phi_inc_i_19(\phi_inc_i[19]~input_o ),
	.phi_inc_i_18(\phi_inc_i[18]~input_o ),
	.phi_inc_i_17(\phi_inc_i[17]~input_o ),
	.phi_inc_i_16(\phi_inc_i[16]~input_o ),
	.phi_inc_i_15(\phi_inc_i[15]~input_o ),
	.phi_inc_i_14(\phi_inc_i[14]~input_o ),
	.phi_inc_i_13(\phi_inc_i[13]~input_o ),
	.phi_inc_i_12(\phi_inc_i[12]~input_o ),
	.phi_inc_i_11(\phi_inc_i[11]~input_o ),
	.phi_inc_i_10(\phi_inc_i[10]~input_o ),
	.phi_inc_i_9(\phi_inc_i[9]~input_o ),
	.phi_inc_i_8(\phi_inc_i[8]~input_o ),
	.phi_inc_i_7(\phi_inc_i[7]~input_o ),
	.phi_inc_i_6(\phi_inc_i[6]~input_o ),
	.phi_inc_i_5(\phi_inc_i[5]~input_o ),
	.phi_inc_i_4(\phi_inc_i[4]~input_o ),
	.phi_inc_i_3(\phi_inc_i[3]~input_o ),
	.phi_inc_i_2(\phi_inc_i[2]~input_o ),
	.phi_inc_i_1(\phi_inc_i[1]~input_o ),
	.phi_inc_i_0(\phi_inc_i[0]~input_o ));

assign \clk~input_o  = clk;

assign \reset_n~input_o  = reset_n;

assign \clken~input_o  = clken;

assign \phi_inc_i[30]~input_o  = phi_inc_i[30];

assign \phi_inc_i[31]~input_o  = phi_inc_i[31];

assign \phi_inc_i[29]~input_o  = phi_inc_i[29];

assign \phi_inc_i[28]~input_o  = phi_inc_i[28];

assign \phi_inc_i[27]~input_o  = phi_inc_i[27];

assign \phi_inc_i[26]~input_o  = phi_inc_i[26];

assign \phi_inc_i[25]~input_o  = phi_inc_i[25];

assign \phi_inc_i[24]~input_o  = phi_inc_i[24];

assign \phi_inc_i[23]~input_o  = phi_inc_i[23];

assign \phi_inc_i[22]~input_o  = phi_inc_i[22];

assign \phi_inc_i[21]~input_o  = phi_inc_i[21];

assign \phi_inc_i[20]~input_o  = phi_inc_i[20];

assign \phi_inc_i[19]~input_o  = phi_inc_i[19];

assign \phi_inc_i[18]~input_o  = phi_inc_i[18];

assign \phi_inc_i[17]~input_o  = phi_inc_i[17];

assign \phi_inc_i[16]~input_o  = phi_inc_i[16];

assign \phi_inc_i[15]~input_o  = phi_inc_i[15];

assign \phi_inc_i[14]~input_o  = phi_inc_i[14];

assign \phi_inc_i[13]~input_o  = phi_inc_i[13];

assign \phi_inc_i[12]~input_o  = phi_inc_i[12];

assign \phi_inc_i[11]~input_o  = phi_inc_i[11];

assign \phi_inc_i[10]~input_o  = phi_inc_i[10];

assign \phi_inc_i[9]~input_o  = phi_inc_i[9];

assign \phi_inc_i[8]~input_o  = phi_inc_i[8];

assign \phi_inc_i[7]~input_o  = phi_inc_i[7];

assign \phi_inc_i[6]~input_o  = phi_inc_i[6];

assign \phi_inc_i[5]~input_o  = phi_inc_i[5];

assign \phi_inc_i[4]~input_o  = phi_inc_i[4];

assign \phi_inc_i[3]~input_o  = phi_inc_i[3];

assign \phi_inc_i[2]~input_o  = phi_inc_i[2];

assign \phi_inc_i[1]~input_o  = phi_inc_i[1];

assign \phi_inc_i[0]~input_o  = phi_inc_i[0];

assign fsin_o[0] = \nco_ii_0|sop|sin_o[0]~q ;

assign fsin_o[1] = \nco_ii_0|sop|sin_o[1]~q ;

assign fsin_o[2] = \nco_ii_0|sop|sin_o[2]~q ;

assign fsin_o[3] = \nco_ii_0|sop|sin_o[3]~q ;

assign fsin_o[4] = \nco_ii_0|sop|sin_o[4]~q ;

assign fsin_o[5] = \nco_ii_0|sop|sin_o[5]~q ;

assign fsin_o[6] = \nco_ii_0|sop|sin_o[6]~q ;

assign fsin_o[7] = \nco_ii_0|sop|sin_o[7]~q ;

assign fsin_o[8] = \nco_ii_0|sop|sin_o[8]~q ;

assign fsin_o[9] = \nco_ii_0|sop|sin_o[9]~q ;

assign fsin_o[10] = \nco_ii_0|sop|sin_o[10]~q ;

assign fsin_o[11] = \nco_ii_0|sop|sin_o[11]~q ;

assign out_valid = \nco_ii_0|ux710isdr|data_ready~q ;

endmodule

module NCO_Lab3_NCO_Lab3_nco_ii_0 (
	sin_o_0,
	sin_o_1,
	sin_o_2,
	sin_o_3,
	sin_o_4,
	sin_o_5,
	sin_o_6,
	sin_o_7,
	sin_o_8,
	sin_o_9,
	sin_o_10,
	sin_o_11,
	data_ready,
	clk,
	reset_n,
	clken,
	phi_inc_i_30,
	phi_inc_i_31,
	phi_inc_i_29,
	phi_inc_i_28,
	phi_inc_i_27,
	phi_inc_i_26,
	phi_inc_i_25,
	phi_inc_i_24,
	phi_inc_i_23,
	phi_inc_i_22,
	phi_inc_i_21,
	phi_inc_i_20,
	phi_inc_i_19,
	phi_inc_i_18,
	phi_inc_i_17,
	phi_inc_i_16,
	phi_inc_i_15,
	phi_inc_i_14,
	phi_inc_i_13,
	phi_inc_i_12,
	phi_inc_i_11,
	phi_inc_i_10,
	phi_inc_i_9,
	phi_inc_i_8,
	phi_inc_i_7,
	phi_inc_i_6,
	phi_inc_i_5,
	phi_inc_i_4,
	phi_inc_i_3,
	phi_inc_i_2,
	phi_inc_i_1,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	sin_o_0;
output 	sin_o_1;
output 	sin_o_2;
output 	sin_o_3;
output 	sin_o_4;
output 	sin_o_5;
output 	sin_o_6;
output 	sin_o_7;
output 	sin_o_8;
output 	sin_o_9;
output 	sin_o_10;
output 	sin_o_11;
output 	data_ready;
input 	clk;
input 	reset_n;
input 	clken;
input 	phi_inc_i_30;
input 	phi_inc_i_31;
input 	phi_inc_i_29;
input 	phi_inc_i_28;
input 	phi_inc_i_27;
input 	phi_inc_i_26;
input 	phi_inc_i_25;
input 	phi_inc_i_24;
input 	phi_inc_i_23;
input 	phi_inc_i_22;
input 	phi_inc_i_21;
input 	phi_inc_i_20;
input 	phi_inc_i_19;
input 	phi_inc_i_18;
input 	phi_inc_i_17;
input 	phi_inc_i_16;
input 	phi_inc_i_15;
input 	phi_inc_i_14;
input 	phi_inc_i_13;
input 	phi_inc_i_12;
input 	phi_inc_i_11;
input 	phi_inc_i_10;
input 	phi_inc_i_9;
input 	phi_inc_i_8;
input 	phi_inc_i_7;
input 	phi_inc_i_6;
input 	phi_inc_i_5;
input 	phi_inc_i_4;
input 	phi_inc_i_3;
input 	phi_inc_i_2;
input 	phi_inc_i_1;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ux002|dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1~portbdataout ;
wire \ux002|dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ;
wire \ux006|sin_o[0]~q ;
wire \ux006|sin_o[1]~q ;
wire \ux006|sin_o[2]~q ;
wire \ux006|sin_o[3]~q ;
wire \ux006|sin_o[4]~q ;
wire \ux006|sin_o[5]~q ;
wire \ux006|sin_o[6]~q ;
wire \ux006|sin_o[7]~q ;
wire \ux006|sin_o[8]~q ;
wire \ux006|sin_o[9]~q ;
wire \ux006|sin_o[10]~q ;
wire \ux006|sin_o[11]~q ;
wire \cordinv|cordic_x_res_2c[0]~q ;
wire \cordinv|cordic_y_res_2c[0]~q ;
wire \cordinv|cordic_y_res_d[1]~q ;
wire \cordinv|cordic_x_res_d[1]~q ;
wire \cordinv|cordic_y_res_2c[1]~q ;
wire \cordinv|cordic_x_res_2c[1]~q ;
wire \cordinv|cordic_y_res_d[2]~q ;
wire \cordinv|cordic_x_res_d[2]~q ;
wire \cordinv|cordic_y_res_2c[2]~q ;
wire \cordinv|cordic_x_res_2c[2]~q ;
wire \cordinv|cordic_y_res_d[3]~q ;
wire \cordinv|cordic_x_res_d[3]~q ;
wire \cordinv|cordic_y_res_2c[3]~q ;
wire \cordinv|cordic_x_res_2c[3]~q ;
wire \cordinv|cordic_y_res_d[4]~q ;
wire \cordinv|cordic_x_res_d[4]~q ;
wire \cordinv|cordic_y_res_2c[4]~q ;
wire \cordinv|cordic_x_res_2c[4]~q ;
wire \cordinv|cordic_y_res_d[5]~q ;
wire \cordinv|cordic_x_res_d[5]~q ;
wire \cordinv|cordic_y_res_2c[5]~q ;
wire \cordinv|cordic_x_res_2c[5]~q ;
wire \cordinv|cordic_y_res_d[6]~q ;
wire \cordinv|cordic_x_res_d[6]~q ;
wire \cordinv|cordic_y_res_2c[6]~q ;
wire \cordinv|cordic_x_res_2c[6]~q ;
wire \cordinv|cordic_y_res_d[7]~q ;
wire \cordinv|cordic_x_res_d[7]~q ;
wire \cordinv|cordic_y_res_2c[7]~q ;
wire \cordinv|cordic_x_res_2c[7]~q ;
wire \cordinv|cordic_y_res_d[8]~q ;
wire \cordinv|cordic_x_res_d[8]~q ;
wire \cordinv|cordic_y_res_2c[8]~q ;
wire \cordinv|cordic_x_res_2c[8]~q ;
wire \cordinv|cordic_y_res_d[9]~q ;
wire \cordinv|cordic_x_res_d[9]~q ;
wire \cordinv|cordic_y_res_2c[9]~q ;
wire \cordinv|cordic_x_res_2c[9]~q ;
wire \cordinv|cordic_y_res_d[10]~q ;
wire \cordinv|cordic_x_res_d[10]~q ;
wire \cordinv|cordic_y_res_2c[10]~q ;
wire \cordinv|cordic_x_res_2c[10]~q ;
wire \cordinv|cordic_y_res_d[11]~q ;
wire \cordinv|cordic_x_res_d[11]~q ;
wire \cordinv|cordic_y_res_2c[11]~q ;
wire \cordinv|cordic_x_res_2c[11]~q ;
wire \u34|u0|auto_generated|dffe1~q ;
wire \u35|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u35|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u34|u0|auto_generated|dffe2~q ;
wire \u35|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u34|u0|auto_generated|dffe3~q ;
wire \u35|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u34|u0|auto_generated|dffe4~q ;
wire \u35|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u34|u0|auto_generated|dffe5~q ;
wire \u35|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u34|u0|auto_generated|dffe6~q ;
wire \u35|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u34|u0|auto_generated|dffe7~q ;
wire \u35|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u34|u0|auto_generated|dffe8~q ;
wire \u35|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u34|u0|auto_generated|dffe9~q ;
wire \u35|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u34|u0|auto_generated|dffe10~q ;
wire \u35|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u34|u0|auto_generated|dffe11~q ;
wire \u35|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u34|u0|auto_generated|dffe12~q ;
wire \ux001|dxxrv[3]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[30]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[31]~q ;
wire \u33|u0|auto_generated|dffe16~q ;
wire \u32|u0|auto_generated|pipeline_dffe[11]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[29]~q ;
wire \u31|u0|auto_generated|dffe12~q ;
wire \u31|u0|auto_generated|dffe1~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[28]~q ;
wire \u32|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u32|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u31|u0|auto_generated|dffe2~q ;
wire \u32|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u31|u0|auto_generated|dffe3~q ;
wire \u32|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u31|u0|auto_generated|dffe4~q ;
wire \u32|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u31|u0|auto_generated|dffe5~q ;
wire \u32|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u31|u0|auto_generated|dffe6~q ;
wire \u32|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u31|u0|auto_generated|dffe7~q ;
wire \u32|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u31|u0|auto_generated|dffe8~q ;
wire \u32|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u31|u0|auto_generated|dffe9~q ;
wire \u32|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u31|u0|auto_generated|dffe10~q ;
wire \u32|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u31|u0|auto_generated|dffe11~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[27]~q ;
wire \u30|u0|auto_generated|dffe16~q ;
wire \u28|u0|auto_generated|dffe12~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[26]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[10]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[25]~q ;
wire \u28|u0|auto_generated|dffe11~q ;
wire \u28|u0|auto_generated|dffe1~q ;
wire \u30|u0|auto_generated|dffe15~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[24]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u28|u0|auto_generated|dffe2~q ;
wire \u29|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u28|u0|auto_generated|dffe3~q ;
wire \u29|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u28|u0|auto_generated|dffe4~q ;
wire \u29|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u28|u0|auto_generated|dffe5~q ;
wire \u29|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u28|u0|auto_generated|dffe6~q ;
wire \u29|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u28|u0|auto_generated|dffe7~q ;
wire \u29|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u28|u0|auto_generated|dffe8~q ;
wire \u29|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u28|u0|auto_generated|dffe9~q ;
wire \u29|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u28|u0|auto_generated|dffe10~q ;
wire \u30|u0|auto_generated|dffe14~q ;
wire \u27|u0|auto_generated|dffe16~q ;
wire \u26|u0|auto_generated|pipeline_dffe[11]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[23]~q ;
wire \u25|u0|auto_generated|dffe12~q ;
wire \u30|u0|auto_generated|dffe13~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[22]~q ;
wire \u26|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u26|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u30|u0|auto_generated|dffe12~q ;
wire \u27|u0|auto_generated|dffe15~q ;
wire \u25|u0|auto_generated|dffe11~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[21]~q ;
wire \u25|u0|auto_generated|dffe10~q ;
wire \u25|u0|auto_generated|dffe1~q ;
wire \u30|u0|auto_generated|dffe11~q ;
wire \u27|u0|auto_generated|dffe14~q ;
wire \u24|u0|auto_generated|dffe16~q ;
wire \u22|u0|auto_generated|dffe12~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[20]~q ;
wire \u23|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u26|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u26|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u25|u0|auto_generated|dffe2~q ;
wire \u26|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u25|u0|auto_generated|dffe3~q ;
wire \u26|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u25|u0|auto_generated|dffe4~q ;
wire \u26|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u25|u0|auto_generated|dffe5~q ;
wire \u26|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u25|u0|auto_generated|dffe6~q ;
wire \u26|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u25|u0|auto_generated|dffe7~q ;
wire \u26|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u25|u0|auto_generated|dffe8~q ;
wire \u26|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u25|u0|auto_generated|dffe9~q ;
wire \u30|u0|auto_generated|dffe10~q ;
wire \u27|u0|auto_generated|dffe13~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[19]~q ;
wire \u30|u0|auto_generated|dffe9~q ;
wire \u27|u0|auto_generated|dffe12~q ;
wire \u24|u0|auto_generated|dffe15~q ;
wire \u23|u0|auto_generated|pipeline_dffe[10]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[18]~q ;
wire \u22|u0|auto_generated|dffe11~q ;
wire \u23|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u23|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u30|u0|auto_generated|dffe8~q ;
wire \u27|u0|auto_generated|dffe11~q ;
wire \u24|u0|auto_generated|dffe14~q ;
wire \u21|u0|auto_generated|dffe16~q ;
wire \u20|u0|auto_generated|pipeline_dffe[11]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[17]~q ;
wire \u22|u0|auto_generated|dffe10~q ;
wire \u19|u0|auto_generated|dffe12~q ;
wire \u22|u0|auto_generated|dffe9~q ;
wire \u22|u0|auto_generated|dffe1~q ;
wire \u30|u0|auto_generated|dffe7~q ;
wire \u27|u0|auto_generated|dffe10~q ;
wire \u24|u0|auto_generated|dffe13~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[16]~q ;
wire \u23|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u23|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u22|u0|auto_generated|dffe2~q ;
wire \u23|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u22|u0|auto_generated|dffe3~q ;
wire \u23|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u22|u0|auto_generated|dffe4~q ;
wire \u23|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u22|u0|auto_generated|dffe5~q ;
wire \u23|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u22|u0|auto_generated|dffe6~q ;
wire \u23|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u22|u0|auto_generated|dffe7~q ;
wire \u23|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u22|u0|auto_generated|dffe8~q ;
wire \u30|u0|auto_generated|dffe6~q ;
wire \u27|u0|auto_generated|dffe9~q ;
wire \u24|u0|auto_generated|dffe12~q ;
wire \u21|u0|auto_generated|dffe15~q ;
wire \u19|u0|auto_generated|dffe11~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[15]~q ;
wire \u20|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u30|u0|auto_generated|dffe5~q ;
wire \u27|u0|auto_generated|dffe8~q ;
wire \u24|u0|auto_generated|dffe11~q ;
wire \u21|u0|auto_generated|dffe14~q ;
wire \u18|u0|auto_generated|dffe16~q ;
wire \u19|u0|auto_generated|dffe10~q ;
wire \u16|u0|auto_generated|dffe12~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[14]~q ;
wire \u20|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u17|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u20|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u20|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u30|u0|auto_generated|dffe4~q ;
wire \u27|u0|auto_generated|dffe7~q ;
wire \u24|u0|auto_generated|dffe10~q ;
wire \u21|u0|auto_generated|dffe13~q ;
wire \u19|u0|auto_generated|dffe9~q ;
wire \ux001|dxxrv[2]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[13]~q ;
wire \u19|u0|auto_generated|dffe8~q ;
wire \u19|u0|auto_generated|dffe1~q ;
wire \u30|u0|auto_generated|dffe3~q ;
wire \u27|u0|auto_generated|dffe6~q ;
wire \u24|u0|auto_generated|dffe9~q ;
wire \u21|u0|auto_generated|dffe12~q ;
wire \u18|u0|auto_generated|dffe15~q ;
wire \u17|u0|auto_generated|pipeline_dffe[10]~q ;
wire \ux001|dxxrv[1]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[12]~q ;
wire \u16|u0|auto_generated|dffe11~q ;
wire \u20|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u20|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u19|u0|auto_generated|dffe2~q ;
wire \u20|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u19|u0|auto_generated|dffe3~q ;
wire \u20|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u19|u0|auto_generated|dffe4~q ;
wire \u20|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u19|u0|auto_generated|dffe5~q ;
wire \u20|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u19|u0|auto_generated|dffe6~q ;
wire \u20|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u19|u0|auto_generated|dffe7~q ;
wire \u30|u0|auto_generated|dffe2~q ;
wire \u27|u0|auto_generated|dffe5~q ;
wire \u24|u0|auto_generated|dffe8~q ;
wire \u21|u0|auto_generated|dffe11~q ;
wire \u18|u0|auto_generated|dffe14~q ;
wire \u15|u0|auto_generated|dffe16~q ;
wire \u17|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u14|u0|auto_generated|pipeline_dffe[11]~q ;
wire \ux001|dxxrv[0]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[11]~q ;
wire \u16|u0|auto_generated|dffe10~q ;
wire \u13|u0|auto_generated|dffe12~q ;
wire \u30|u0|auto_generated|dffe1~q ;
wire \u27|u0|auto_generated|dffe4~q ;
wire \u24|u0|auto_generated|dffe7~q ;
wire \u21|u0|auto_generated|dffe10~q ;
wire \u18|u0|auto_generated|dffe13~q ;
wire \u17|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u16|u0|auto_generated|dffe9~q ;
wire \u17|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u17|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u27|u0|auto_generated|dffe3~q ;
wire \u24|u0|auto_generated|dffe6~q ;
wire \u21|u0|auto_generated|dffe9~q ;
wire \u18|u0|auto_generated|dffe12~q ;
wire \u15|u0|auto_generated|dffe15~q ;
wire \u13|u0|auto_generated|dffe11~q ;
wire \u16|u0|auto_generated|dffe8~q ;
wire \u14|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u16|u0|auto_generated|dffe7~q ;
wire \u16|u0|auto_generated|dffe1~q ;
wire \u27|u0|auto_generated|dffe2~q ;
wire \u24|u0|auto_generated|dffe5~q ;
wire \u21|u0|auto_generated|dffe8~q ;
wire \u18|u0|auto_generated|dffe11~q ;
wire \u15|u0|auto_generated|dffe14~q ;
wire \u12|u0|auto_generated|dffe16~q ;
wire \u13|u0|auto_generated|dffe10~q ;
wire \u10|u0|auto_generated|dffe12~q ;
wire \u14|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u11|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u17|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u17|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u16|u0|auto_generated|dffe2~q ;
wire \u17|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u16|u0|auto_generated|dffe3~q ;
wire \u17|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u16|u0|auto_generated|dffe4~q ;
wire \u17|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u16|u0|auto_generated|dffe5~q ;
wire \u17|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u16|u0|auto_generated|dffe6~q ;
wire \u27|u0|auto_generated|dffe1~q ;
wire \u24|u0|auto_generated|dffe4~q ;
wire \u21|u0|auto_generated|dffe7~q ;
wire \u18|u0|auto_generated|dffe10~q ;
wire \u15|u0|auto_generated|dffe13~q ;
wire \u13|u0|auto_generated|dffe9~q ;
wire \u14|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u24|u0|auto_generated|dffe3~q ;
wire \u21|u0|auto_generated|dffe6~q ;
wire \u18|u0|auto_generated|dffe9~q ;
wire \u15|u0|auto_generated|dffe12~q ;
wire \u12|u0|auto_generated|dffe15~q ;
wire \u13|u0|auto_generated|dffe8~q ;
wire \u11|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u14|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u10|u0|auto_generated|dffe11~q ;
wire \u14|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u14|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u24|u0|auto_generated|dffe2~q ;
wire \u21|u0|auto_generated|dffe5~q ;
wire \u18|u0|auto_generated|dffe8~q ;
wire \u15|u0|auto_generated|dffe11~q ;
wire \u12|u0|auto_generated|dffe14~q ;
wire \u9|u0|auto_generated|dffe16~q ;
wire \u13|u0|auto_generated|dffe7~q ;
wire \u11|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u8|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u10|u0|auto_generated|dffe10~q ;
wire \u7|u0|auto_generated|dffe12~q ;
wire \u13|u0|auto_generated|dffe6~q ;
wire \u13|u0|auto_generated|dffe1~q ;
wire \u24|u0|auto_generated|dffe1~q ;
wire \u21|u0|auto_generated|dffe4~q ;
wire \u18|u0|auto_generated|dffe7~q ;
wire \u15|u0|auto_generated|dffe10~q ;
wire \u12|u0|auto_generated|dffe13~q ;
wire \u11|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u10|u0|auto_generated|dffe9~q ;
wire \u14|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u14|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u13|u0|auto_generated|dffe2~q ;
wire \u14|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u13|u0|auto_generated|dffe3~q ;
wire \u14|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u13|u0|auto_generated|dffe4~q ;
wire \u14|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u13|u0|auto_generated|dffe5~q ;
wire \u21|u0|auto_generated|dffe3~q ;
wire \u18|u0|auto_generated|dffe6~q ;
wire \u15|u0|auto_generated|dffe9~q ;
wire \u12|u0|auto_generated|dffe12~q ;
wire \u9|u0|auto_generated|dffe15~q ;
wire \u8|a[0]~q ;
wire \u11|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u7|u0|auto_generated|dffe11~q ;
wire \u10|u0|auto_generated|dffe8~q ;
wire \u8|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u21|u0|auto_generated|dffe2~q ;
wire \u18|u0|auto_generated|dffe5~q ;
wire \u15|u0|auto_generated|dffe8~q ;
wire \u12|u0|auto_generated|dffe11~q ;
wire \u9|u0|auto_generated|dffe14~q ;
wire \u6|u0|auto_generated|dffe16~q ;
wire \u11|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u7|u0|auto_generated|dffe10~q ;
wire \u5|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u4|u0|auto_generated|dffe12~q ;
wire \u10|u0|auto_generated|dffe7~q ;
wire \u8|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u11|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u11|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u21|u0|auto_generated|dffe1~q ;
wire \u18|u0|auto_generated|dffe4~q ;
wire \u15|u0|auto_generated|dffe7~q ;
wire \u12|u0|auto_generated|dffe10~q ;
wire \u9|u0|auto_generated|dffe13~q ;
wire \u7|u0|auto_generated|dffe9~q ;
wire \u5|a[0]~q ;
wire \u5|xordvalue[2]~q ;
wire \u5|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u10|u0|auto_generated|dffe6~q ;
wire \u8|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u10|u0|auto_generated|dffe5~q ;
wire \u10|u0|auto_generated|dffe1~q ;
wire \u18|u0|auto_generated|dffe3~q ;
wire \u15|u0|auto_generated|dffe6~q ;
wire \u12|u0|auto_generated|dffe9~q ;
wire \u9|u0|auto_generated|dffe12~q ;
wire \u6|u0|auto_generated|dffe15~q ;
wire \u7|u0|auto_generated|dffe8~q ;
wire \u3|u0|auto_generated|dffe16~q ;
wire \cfs|cor1x[10]~q ;
wire \u5|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u8|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u4|u0|auto_generated|dffe11~q ;
wire \u11|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u11|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u10|u0|auto_generated|dffe2~q ;
wire \u11|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u10|u0|auto_generated|dffe3~q ;
wire \u11|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u10|u0|auto_generated|dffe4~q ;
wire \u18|u0|auto_generated|dffe2~q ;
wire \u15|u0|auto_generated|dffe5~q ;
wire \u12|u0|auto_generated|dffe8~q ;
wire \u9|u0|auto_generated|dffe11~q ;
wire \u6|u0|auto_generated|dffe14~q ;
wire \u7|u0|auto_generated|dffe7~q ;
wire \ci|corx[10]~q ;
wire \u5|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u8|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u4|u0|auto_generated|dffe10~q ;
wire \u18|u0|auto_generated|dffe1~q ;
wire \u15|u0|auto_generated|dffe4~q ;
wire \u12|u0|auto_generated|dffe7~q ;
wire \u9|u0|auto_generated|dffe10~q ;
wire \u6|u0|auto_generated|dffe13~q ;
wire \u7|u0|auto_generated|dffe6~q ;
wire \u5|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u8|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u4|u0|auto_generated|dffe9~q ;
wire \u8|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u8|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u15|u0|auto_generated|dffe3~q ;
wire \u12|u0|auto_generated|dffe6~q ;
wire \u9|u0|auto_generated|dffe9~q ;
wire \u6|u0|auto_generated|dffe12~q ;
wire \u3|u0|auto_generated|dffe15~q ;
wire \u7|u0|auto_generated|dffe5~q ;
wire \u5|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u4|u0|auto_generated|dffe8~q ;
wire \u7|u0|auto_generated|dffe4~q ;
wire \u7|u0|auto_generated|dffe1~q ;
wire \u15|u0|auto_generated|dffe2~q ;
wire \u12|u0|auto_generated|dffe5~q ;
wire \u9|u0|auto_generated|dffe8~q ;
wire \u6|u0|auto_generated|dffe11~q ;
wire \u3|u0|auto_generated|dffe14~q ;
wire \ci|corz[14]~q ;
wire \u5|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u4|u0|auto_generated|dffe7~q ;
wire \u8|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u8|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u7|u0|auto_generated|dffe2~q ;
wire \u8|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u7|u0|auto_generated|dffe3~q ;
wire \u15|u0|auto_generated|dffe1~q ;
wire \u12|u0|auto_generated|dffe4~q ;
wire \u9|u0|auto_generated|dffe7~q ;
wire \u6|u0|auto_generated|dffe10~q ;
wire \u3|u0|auto_generated|dffe13~q ;
wire \ux002|dxxpdo[18]~q ;
wire \ci|corz[13]~q ;
wire \u5|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u4|u0|auto_generated|dffe6~q ;
wire \u5|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u12|u0|auto_generated|dffe3~q ;
wire \u9|u0|auto_generated|dffe6~q ;
wire \u6|u0|auto_generated|dffe9~q ;
wire \u3|u0|auto_generated|dffe12~q ;
wire \ux002|dxxpdo[17]~q ;
wire \ci|corz[12]~q ;
wire \u4|u0|auto_generated|dffe5~q ;
wire \u5|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u12|u0|auto_generated|dffe2~q ;
wire \u9|u0|auto_generated|dffe5~q ;
wire \u6|u0|auto_generated|dffe8~q ;
wire \u3|u0|auto_generated|dffe11~q ;
wire \ux002|dxxpdo[16]~q ;
wire \ci|corz[11]~q ;
wire \u4|u0|auto_generated|dffe4~q ;
wire \u4|u0|auto_generated|dffe3~q ;
wire \u4|u0|auto_generated|dffe1~q ;
wire \u12|u0|auto_generated|dffe1~q ;
wire \u9|u0|auto_generated|dffe4~q ;
wire \u6|u0|auto_generated|dffe7~q ;
wire \u3|u0|auto_generated|dffe10~q ;
wire \ux002|dxxpdo[15]~q ;
wire \ci|corz[10]~q ;
wire \u4|u0|auto_generated|dffe2~q ;
wire \u9|u0|auto_generated|dffe3~q ;
wire \u6|u0|auto_generated|dffe6~q ;
wire \u3|u0|auto_generated|dffe9~q ;
wire \ux002|dxxpdo[14]~q ;
wire \ci|corz[9]~q ;
wire \u9|u0|auto_generated|dffe2~q ;
wire \u6|u0|auto_generated|dffe5~q ;
wire \u3|u0|auto_generated|dffe8~q ;
wire \ux002|dxxpdo[13]~q ;
wire \ci|corz[8]~q ;
wire \u9|u0|auto_generated|dffe1~q ;
wire \u6|u0|auto_generated|dffe4~q ;
wire \u3|u0|auto_generated|dffe7~q ;
wire \ux002|dxxpdo[12]~q ;
wire \ci|corz[7]~q ;
wire \u6|u0|auto_generated|dffe3~q ;
wire \u3|u0|auto_generated|dffe6~q ;
wire \ux002|dxxpdo[11]~q ;
wire \ci|corz[6]~q ;
wire \u6|u0|auto_generated|dffe2~q ;
wire \u3|u0|auto_generated|dffe5~q ;
wire \ux002|dxxpdo[10]~q ;
wire \ci|corz[5]~q ;
wire \u6|u0|auto_generated|dffe1~q ;
wire \u3|u0|auto_generated|dffe4~q ;
wire \ux002|dxxpdo[9]~q ;
wire \ci|corz[4]~q ;
wire \u3|u0|auto_generated|dffe3~q ;
wire \ux002|dxxpdo[8]~q ;
wire \ci|corz[3]~q ;
wire \u3|u0|auto_generated|dffe2~q ;
wire \ux002|dxxpdo[7]~q ;
wire \ci|corz[2]~q ;
wire \u3|u0|auto_generated|dffe1~q ;
wire \ux002|dxxpdo[6]~q ;
wire \ci|corz[1]~q ;
wire \ux002|dxxpdo[5]~q ;
wire \ci|corz[0]~q ;
wire \ux002|dxxpdo[4]~q ;


NCO_Lab3_cordic_zxor_1p_lpm_10 u9(
	.dffe16(\u9|u0|auto_generated|dffe16~q ),
	.dffe15(\u9|u0|auto_generated|dffe15~q ),
	.a_0(\u8|a[0]~q ),
	.dffe14(\u9|u0|auto_generated|dffe14~q ),
	.dffe161(\u6|u0|auto_generated|dffe16~q ),
	.dffe13(\u9|u0|auto_generated|dffe13~q ),
	.dffe12(\u9|u0|auto_generated|dffe12~q ),
	.dffe151(\u6|u0|auto_generated|dffe15~q ),
	.dffe11(\u9|u0|auto_generated|dffe11~q ),
	.dffe141(\u6|u0|auto_generated|dffe14~q ),
	.dffe10(\u9|u0|auto_generated|dffe10~q ),
	.dffe131(\u6|u0|auto_generated|dffe13~q ),
	.dffe9(\u9|u0|auto_generated|dffe9~q ),
	.dffe121(\u6|u0|auto_generated|dffe12~q ),
	.dffe8(\u9|u0|auto_generated|dffe8~q ),
	.dffe111(\u6|u0|auto_generated|dffe11~q ),
	.dffe7(\u9|u0|auto_generated|dffe7~q ),
	.dffe101(\u6|u0|auto_generated|dffe10~q ),
	.dffe6(\u9|u0|auto_generated|dffe6~q ),
	.dffe91(\u6|u0|auto_generated|dffe9~q ),
	.dffe5(\u9|u0|auto_generated|dffe5~q ),
	.dffe81(\u6|u0|auto_generated|dffe8~q ),
	.dffe4(\u9|u0|auto_generated|dffe4~q ),
	.dffe71(\u6|u0|auto_generated|dffe7~q ),
	.dffe3(\u9|u0|auto_generated|dffe3~q ),
	.dffe61(\u6|u0|auto_generated|dffe6~q ),
	.dffe2(\u9|u0|auto_generated|dffe2~q ),
	.dffe51(\u6|u0|auto_generated|dffe5~q ),
	.dffe1(\u9|u0|auto_generated|dffe1~q ),
	.dffe41(\u6|u0|auto_generated|dffe4~q ),
	.dffe31(\u6|u0|auto_generated|dffe3~q ),
	.dffe21(\u6|u0|auto_generated|dffe2~q ),
	.dffe17(\u6|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm_10 u8(
	.pipeline_dffe_11(\u8|u0|auto_generated|pipeline_dffe[11]~q ),
	.a_0(\u8|a[0]~q ),
	.pipeline_dffe_10(\u8|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe16(\u6|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_111(\u5|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe12(\u4|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_9(\u8|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\u5|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_8(\u8|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u5|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_7(\u8|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe11(\u4|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_81(\u5|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_6(\u8|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe10(\u4|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_71(\u5|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_5(\u8|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe9(\u4|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_3(\u8|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u8|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_61(\u5|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe8(\u4|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_51(\u5|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe7(\u4|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_0(\u8|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u8|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u8|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_41(\u5|u0|auto_generated|pipeline_dffe[4]~q ),
	.dffe6(\u4|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_31(\u5|u0|auto_generated|pipeline_dffe[3]~q ),
	.dffe5(\u4|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_21(\u5|u0|auto_generated|pipeline_dffe[2]~q ),
	.dffe4(\u4|u0|auto_generated|dffe4~q ),
	.dffe3(\u4|u0|auto_generated|dffe3~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm_10 u7(
	.dffe12(\u7|u0|auto_generated|dffe12~q ),
	.dffe11(\u7|u0|auto_generated|dffe11~q ),
	.dffe16(\u6|u0|auto_generated|dffe16~q ),
	.dffe10(\u7|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_11(\u5|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe121(\u4|u0|auto_generated|dffe12~q ),
	.dffe9(\u7|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_10(\u5|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe8(\u7|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_9(\u5|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe111(\u4|u0|auto_generated|dffe11~q ),
	.dffe7(\u7|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_8(\u5|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe101(\u4|u0|auto_generated|dffe10~q ),
	.dffe6(\u7|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_7(\u5|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe91(\u4|u0|auto_generated|dffe9~q ),
	.dffe5(\u7|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_6(\u5|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe81(\u4|u0|auto_generated|dffe8~q ),
	.dffe4(\u7|u0|auto_generated|dffe4~q ),
	.dffe1(\u7|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_5(\u5|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe71(\u4|u0|auto_generated|dffe7~q ),
	.dffe2(\u7|u0|auto_generated|dffe2~q ),
	.dffe3(\u7|u0|auto_generated|dffe3~q ),
	.pipeline_dffe_4(\u5|u0|auto_generated|pipeline_dffe[4]~q ),
	.dffe61(\u4|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_3(\u5|u0|auto_generated|pipeline_dffe[3]~q ),
	.dffe51(\u4|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_2(\u5|u0|auto_generated|pipeline_dffe[2]~q ),
	.dffe41(\u4|u0|auto_generated|dffe4~q ),
	.dffe31(\u4|u0|auto_generated|dffe3~q ),
	.dffe13(\u4|u0|auto_generated|dffe1~q ),
	.dffe21(\u4|u0|auto_generated|dffe2~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_zxor_1p_lpm_9 u6(
	.dffe16(\u6|u0|auto_generated|dffe16~q ),
	.a_0(\u5|a[0]~q ),
	.dffe15(\u6|u0|auto_generated|dffe15~q ),
	.dffe161(\u3|u0|auto_generated|dffe16~q ),
	.dffe14(\u6|u0|auto_generated|dffe14~q ),
	.dffe13(\u6|u0|auto_generated|dffe13~q ),
	.dffe12(\u6|u0|auto_generated|dffe12~q ),
	.dffe151(\u3|u0|auto_generated|dffe15~q ),
	.dffe11(\u6|u0|auto_generated|dffe11~q ),
	.dffe141(\u3|u0|auto_generated|dffe14~q ),
	.dffe10(\u6|u0|auto_generated|dffe10~q ),
	.dffe131(\u3|u0|auto_generated|dffe13~q ),
	.dffe9(\u6|u0|auto_generated|dffe9~q ),
	.dffe121(\u3|u0|auto_generated|dffe12~q ),
	.dffe8(\u6|u0|auto_generated|dffe8~q ),
	.dffe111(\u3|u0|auto_generated|dffe11~q ),
	.dffe7(\u6|u0|auto_generated|dffe7~q ),
	.dffe101(\u3|u0|auto_generated|dffe10~q ),
	.dffe6(\u6|u0|auto_generated|dffe6~q ),
	.dffe91(\u3|u0|auto_generated|dffe9~q ),
	.dffe5(\u6|u0|auto_generated|dffe5~q ),
	.dffe81(\u3|u0|auto_generated|dffe8~q ),
	.dffe4(\u6|u0|auto_generated|dffe4~q ),
	.dffe71(\u3|u0|auto_generated|dffe7~q ),
	.dffe3(\u6|u0|auto_generated|dffe3~q ),
	.dffe61(\u3|u0|auto_generated|dffe6~q ),
	.dffe2(\u6|u0|auto_generated|dffe2~q ),
	.dffe51(\u3|u0|auto_generated|dffe5~q ),
	.dffe1(\u6|u0|auto_generated|dffe1~q ),
	.dffe41(\u3|u0|auto_generated|dffe4~q ),
	.dffe31(\u3|u0|auto_generated|dffe3~q ),
	.dffe21(\u3|u0|auto_generated|dffe2~q ),
	.dffe17(\u3|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm_9 u5(
	.pipeline_dffe_11(\u5|u0|auto_generated|pipeline_dffe[11]~q ),
	.a_0(\u5|a[0]~q ),
	.xordvalue_2(\u5|xordvalue[2]~q ),
	.pipeline_dffe_10(\u5|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe16(\u3|u0|auto_generated|dffe16~q ),
	.cor1x_10(\cfs|cor1x[10]~q ),
	.pipeline_dffe_9(\u5|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\u5|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\u5|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\u5|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\u5|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\u5|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\u5|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\u5|u0|auto_generated|pipeline_dffe[2]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm_9 u4(
	.dffe12(\u4|u0|auto_generated|dffe12~q ),
	.a_0(\u5|a[0]~q ),
	.xordvalue_2(\u5|xordvalue[2]~q ),
	.dffe16(\u3|u0|auto_generated|dffe16~q ),
	.cor1x_10(\cfs|cor1x[10]~q ),
	.dffe11(\u4|u0|auto_generated|dffe11~q ),
	.dffe10(\u4|u0|auto_generated|dffe10~q ),
	.dffe9(\u4|u0|auto_generated|dffe9~q ),
	.dffe8(\u4|u0|auto_generated|dffe8~q ),
	.dffe7(\u4|u0|auto_generated|dffe7~q ),
	.dffe6(\u4|u0|auto_generated|dffe6~q ),
	.dffe5(\u4|u0|auto_generated|dffe5~q ),
	.dffe4(\u4|u0|auto_generated|dffe4~q ),
	.dffe3(\u4|u0|auto_generated|dffe3~q ),
	.dffe1(\u4|u0|auto_generated|dffe1~q ),
	.dffe2(\u4|u0|auto_generated|dffe2~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_zxor_1p_lpm_6 u3(
	.dffe16(\u3|u0|auto_generated|dffe16~q ),
	.corx_10(\ci|corx[10]~q ),
	.dffe15(\u3|u0|auto_generated|dffe15~q ),
	.dffe14(\u3|u0|auto_generated|dffe14~q ),
	.corz_14(\ci|corz[14]~q ),
	.dffe13(\u3|u0|auto_generated|dffe13~q ),
	.corz_13(\ci|corz[13]~q ),
	.dffe12(\u3|u0|auto_generated|dffe12~q ),
	.corz_12(\ci|corz[12]~q ),
	.dffe11(\u3|u0|auto_generated|dffe11~q ),
	.corz_11(\ci|corz[11]~q ),
	.dffe10(\u3|u0|auto_generated|dffe10~q ),
	.corz_10(\ci|corz[10]~q ),
	.dffe9(\u3|u0|auto_generated|dffe9~q ),
	.corz_9(\ci|corz[9]~q ),
	.dffe8(\u3|u0|auto_generated|dffe8~q ),
	.corz_8(\ci|corz[8]~q ),
	.dffe7(\u3|u0|auto_generated|dffe7~q ),
	.corz_7(\ci|corz[7]~q ),
	.dffe6(\u3|u0|auto_generated|dffe6~q ),
	.corz_6(\ci|corz[6]~q ),
	.dffe5(\u3|u0|auto_generated|dffe5~q ),
	.corz_5(\ci|corz[5]~q ),
	.dffe4(\u3|u0|auto_generated|dffe4~q ),
	.corz_4(\ci|corz[4]~q ),
	.dffe3(\u3|u0|auto_generated|dffe3~q ),
	.corz_3(\ci|corz[3]~q ),
	.dffe2(\u3|u0|auto_generated|dffe2~q ),
	.corz_2(\ci|corz[2]~q ),
	.dffe1(\u3|u0|auto_generated|dffe1~q ),
	.corz_1(\ci|corz[1]~q ),
	.corz_0(\ci|corz[0]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_asj_dxx ux002(
	.ram_block8a1(\ux002|dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1~portbdataout ),
	.ram_block8a0(\ux002|dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ),
	.dxxrv_3(\ux001|dxxrv[3]~q ),
	.pipeline_dffe_30(\ux000|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_31(\ux000|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_29(\ux000|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_28(\ux000|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_27(\ux000|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_26(\ux000|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_25(\ux000|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_24(\ux000|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_23(\ux000|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_22(\ux000|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_21(\ux000|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_20(\ux000|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_19(\ux000|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_18(\ux000|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_17(\ux000|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\ux000|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_15(\ux000|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_14(\ux000|acc|auto_generated|pipeline_dffe[14]~q ),
	.dxxrv_2(\ux001|dxxrv[2]~q ),
	.pipeline_dffe_13(\ux000|acc|auto_generated|pipeline_dffe[13]~q ),
	.dxxrv_1(\ux001|dxxrv[1]~q ),
	.pipeline_dffe_12(\ux000|acc|auto_generated|pipeline_dffe[12]~q ),
	.dxxrv_0(\ux001|dxxrv[0]~q ),
	.pipeline_dffe_11(\ux000|acc|auto_generated|pipeline_dffe[11]~q ),
	.dxxpdo_18(\ux002|dxxpdo[18]~q ),
	.dxxpdo_17(\ux002|dxxpdo[17]~q ),
	.dxxpdo_16(\ux002|dxxpdo[16]~q ),
	.dxxpdo_15(\ux002|dxxpdo[15]~q ),
	.dxxpdo_14(\ux002|dxxpdo[14]~q ),
	.dxxpdo_13(\ux002|dxxpdo[13]~q ),
	.dxxpdo_12(\ux002|dxxpdo[12]~q ),
	.dxxpdo_11(\ux002|dxxpdo[11]~q ),
	.dxxpdo_10(\ux002|dxxpdo[10]~q ),
	.dxxpdo_9(\ux002|dxxpdo[9]~q ),
	.dxxpdo_8(\ux002|dxxpdo[8]~q ),
	.dxxpdo_7(\ux002|dxxpdo[7]~q ),
	.dxxpdo_6(\ux002|dxxpdo[6]~q ),
	.dxxpdo_5(\ux002|dxxpdo[5]~q ),
	.dxxpdo_4(\ux002|dxxpdo[4]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_asj_dxx_g ux001(
	.dxxrv_3(\ux001|dxxrv[3]~q ),
	.dxxrv_2(\ux001|dxxrv[2]~q ),
	.dxxrv_1(\ux001|dxxrv[1]~q ),
	.dxxrv_0(\ux001|dxxrv[0]~q ),
	.clk(clk),
	.reset(reset_n),
	.clken(clken));

NCO_Lab3_asj_altqmcpipe ux000(
	.pipeline_dffe_30(\ux000|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_31(\ux000|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_29(\ux000|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_28(\ux000|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_27(\ux000|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_26(\ux000|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_25(\ux000|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_24(\ux000|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_23(\ux000|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_22(\ux000|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_21(\ux000|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_20(\ux000|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_19(\ux000|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_18(\ux000|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_17(\ux000|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\ux000|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_15(\ux000|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_14(\ux000|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\ux000|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_12(\ux000|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\ux000|acc|auto_generated|pipeline_dffe[11]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken),
	.phi_inc_i_30(phi_inc_i_30),
	.phi_inc_i_31(phi_inc_i_31),
	.phi_inc_i_29(phi_inc_i_29),
	.phi_inc_i_28(phi_inc_i_28),
	.phi_inc_i_27(phi_inc_i_27),
	.phi_inc_i_26(phi_inc_i_26),
	.phi_inc_i_25(phi_inc_i_25),
	.phi_inc_i_24(phi_inc_i_24),
	.phi_inc_i_23(phi_inc_i_23),
	.phi_inc_i_22(phi_inc_i_22),
	.phi_inc_i_21(phi_inc_i_21),
	.phi_inc_i_20(phi_inc_i_20),
	.phi_inc_i_19(phi_inc_i_19),
	.phi_inc_i_18(phi_inc_i_18),
	.phi_inc_i_17(phi_inc_i_17),
	.phi_inc_i_16(phi_inc_i_16),
	.phi_inc_i_15(phi_inc_i_15),
	.phi_inc_i_14(phi_inc_i_14),
	.phi_inc_i_13(phi_inc_i_13),
	.phi_inc_i_12(phi_inc_i_12),
	.phi_inc_i_11(phi_inc_i_11),
	.phi_inc_i_10(phi_inc_i_10),
	.phi_inc_i_9(phi_inc_i_9),
	.phi_inc_i_8(phi_inc_i_8),
	.phi_inc_i_7(phi_inc_i_7),
	.phi_inc_i_6(phi_inc_i_6),
	.phi_inc_i_5(phi_inc_i_5),
	.phi_inc_i_4(phi_inc_i_4),
	.phi_inc_i_3(phi_inc_i_3),
	.phi_inc_i_2(phi_inc_i_2),
	.phi_inc_i_1(phi_inc_i_1),
	.phi_inc_i_0(phi_inc_i_0));

NCO_Lab3_cord_fs cfs(
	.cor1x_10(\cfs|cor1x[10]~q ),
	.corx_10(\ci|corx[10]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cord_init ci(
	.corx_10(\ci|corx[10]~q ),
	.corz_14(\ci|corz[14]~q ),
	.dxxpdo_18(\ux002|dxxpdo[18]~q ),
	.corz_13(\ci|corz[13]~q ),
	.dxxpdo_17(\ux002|dxxpdo[17]~q ),
	.corz_12(\ci|corz[12]~q ),
	.dxxpdo_16(\ux002|dxxpdo[16]~q ),
	.corz_11(\ci|corz[11]~q ),
	.dxxpdo_15(\ux002|dxxpdo[15]~q ),
	.corz_10(\ci|corz[10]~q ),
	.dxxpdo_14(\ux002|dxxpdo[14]~q ),
	.corz_9(\ci|corz[9]~q ),
	.dxxpdo_13(\ux002|dxxpdo[13]~q ),
	.corz_8(\ci|corz[8]~q ),
	.dxxpdo_12(\ux002|dxxpdo[12]~q ),
	.corz_7(\ci|corz[7]~q ),
	.dxxpdo_11(\ux002|dxxpdo[11]~q ),
	.corz_6(\ci|corz[6]~q ),
	.dxxpdo_10(\ux002|dxxpdo[10]~q ),
	.corz_5(\ci|corz[5]~q ),
	.dxxpdo_9(\ux002|dxxpdo[9]~q ),
	.corz_4(\ci|corz[4]~q ),
	.dxxpdo_8(\ux002|dxxpdo[8]~q ),
	.corz_3(\ci|corz[3]~q ),
	.dxxpdo_7(\ux002|dxxpdo[7]~q ),
	.corz_2(\ci|corz[2]~q ),
	.dxxpdo_6(\ux002|dxxpdo[6]~q ),
	.corz_1(\ci|corz[1]~q ),
	.dxxpdo_5(\ux002|dxxpdo[5]~q ),
	.corz_0(\ci|corz[0]~q ),
	.dxxpdo_4(\ux002|dxxpdo[4]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_sop_reg sop(
	.sin_o_0(sin_o_0),
	.sin_o_1(sin_o_1),
	.sin_o_2(sin_o_2),
	.sin_o_3(sin_o_3),
	.sin_o_4(sin_o_4),
	.sin_o_5(sin_o_5),
	.sin_o_6(sin_o_6),
	.sin_o_7(sin_o_7),
	.sin_o_8(sin_o_8),
	.sin_o_9(sin_o_9),
	.sin_o_10(sin_o_10),
	.sin_o_11(sin_o_11),
	.sin_o_01(\ux006|sin_o[0]~q ),
	.sin_o_12(\ux006|sin_o[1]~q ),
	.sin_o_21(\ux006|sin_o[2]~q ),
	.sin_o_31(\ux006|sin_o[3]~q ),
	.sin_o_41(\ux006|sin_o[4]~q ),
	.sin_o_51(\ux006|sin_o[5]~q ),
	.sin_o_61(\ux006|sin_o[6]~q ),
	.sin_o_71(\ux006|sin_o[7]~q ),
	.sin_o_81(\ux006|sin_o[8]~q ),
	.sin_o_91(\ux006|sin_o[9]~q ),
	.sin_o_101(\ux006|sin_o[10]~q ),
	.sin_o_111(\ux006|sin_o[11]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_asj_crs_par ux006(
	.ram_block8a1(\ux002|dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1~portbdataout ),
	.ram_block8a0(\ux002|dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0~portbdataout ),
	.sin_o_0(\ux006|sin_o[0]~q ),
	.sin_o_1(\ux006|sin_o[1]~q ),
	.sin_o_2(\ux006|sin_o[2]~q ),
	.sin_o_3(\ux006|sin_o[3]~q ),
	.sin_o_4(\ux006|sin_o[4]~q ),
	.sin_o_5(\ux006|sin_o[5]~q ),
	.sin_o_6(\ux006|sin_o[6]~q ),
	.sin_o_7(\ux006|sin_o[7]~q ),
	.sin_o_8(\ux006|sin_o[8]~q ),
	.sin_o_9(\ux006|sin_o[9]~q ),
	.sin_o_10(\ux006|sin_o[10]~q ),
	.sin_o_11(\ux006|sin_o[11]~q ),
	.cordic_x_res_2c_0(\cordinv|cordic_x_res_2c[0]~q ),
	.cordic_y_res_2c_0(\cordinv|cordic_y_res_2c[0]~q ),
	.cordic_y_res_d_1(\cordinv|cordic_y_res_d[1]~q ),
	.cordic_x_res_d_1(\cordinv|cordic_x_res_d[1]~q ),
	.cordic_y_res_2c_1(\cordinv|cordic_y_res_2c[1]~q ),
	.cordic_x_res_2c_1(\cordinv|cordic_x_res_2c[1]~q ),
	.cordic_y_res_d_2(\cordinv|cordic_y_res_d[2]~q ),
	.cordic_x_res_d_2(\cordinv|cordic_x_res_d[2]~q ),
	.cordic_y_res_2c_2(\cordinv|cordic_y_res_2c[2]~q ),
	.cordic_x_res_2c_2(\cordinv|cordic_x_res_2c[2]~q ),
	.cordic_y_res_d_3(\cordinv|cordic_y_res_d[3]~q ),
	.cordic_x_res_d_3(\cordinv|cordic_x_res_d[3]~q ),
	.cordic_y_res_2c_3(\cordinv|cordic_y_res_2c[3]~q ),
	.cordic_x_res_2c_3(\cordinv|cordic_x_res_2c[3]~q ),
	.cordic_y_res_d_4(\cordinv|cordic_y_res_d[4]~q ),
	.cordic_x_res_d_4(\cordinv|cordic_x_res_d[4]~q ),
	.cordic_y_res_2c_4(\cordinv|cordic_y_res_2c[4]~q ),
	.cordic_x_res_2c_4(\cordinv|cordic_x_res_2c[4]~q ),
	.cordic_y_res_d_5(\cordinv|cordic_y_res_d[5]~q ),
	.cordic_x_res_d_5(\cordinv|cordic_x_res_d[5]~q ),
	.cordic_y_res_2c_5(\cordinv|cordic_y_res_2c[5]~q ),
	.cordic_x_res_2c_5(\cordinv|cordic_x_res_2c[5]~q ),
	.cordic_y_res_d_6(\cordinv|cordic_y_res_d[6]~q ),
	.cordic_x_res_d_6(\cordinv|cordic_x_res_d[6]~q ),
	.cordic_y_res_2c_6(\cordinv|cordic_y_res_2c[6]~q ),
	.cordic_x_res_2c_6(\cordinv|cordic_x_res_2c[6]~q ),
	.cordic_y_res_d_7(\cordinv|cordic_y_res_d[7]~q ),
	.cordic_x_res_d_7(\cordinv|cordic_x_res_d[7]~q ),
	.cordic_y_res_2c_7(\cordinv|cordic_y_res_2c[7]~q ),
	.cordic_x_res_2c_7(\cordinv|cordic_x_res_2c[7]~q ),
	.cordic_y_res_d_8(\cordinv|cordic_y_res_d[8]~q ),
	.cordic_x_res_d_8(\cordinv|cordic_x_res_d[8]~q ),
	.cordic_y_res_2c_8(\cordinv|cordic_y_res_2c[8]~q ),
	.cordic_x_res_2c_8(\cordinv|cordic_x_res_2c[8]~q ),
	.cordic_y_res_d_9(\cordinv|cordic_y_res_d[9]~q ),
	.cordic_x_res_d_9(\cordinv|cordic_x_res_d[9]~q ),
	.cordic_y_res_2c_9(\cordinv|cordic_y_res_2c[9]~q ),
	.cordic_x_res_2c_9(\cordinv|cordic_x_res_2c[9]~q ),
	.cordic_y_res_d_10(\cordinv|cordic_y_res_d[10]~q ),
	.cordic_x_res_d_10(\cordinv|cordic_x_res_d[10]~q ),
	.cordic_y_res_2c_10(\cordinv|cordic_y_res_2c[10]~q ),
	.cordic_x_res_2c_10(\cordinv|cordic_x_res_2c[10]~q ),
	.cordic_y_res_d_11(\cordinv|cordic_y_res_d[11]~q ),
	.cordic_x_res_d_11(\cordinv|cordic_x_res_d[11]~q ),
	.cordic_y_res_2c_11(\cordinv|cordic_y_res_2c[11]~q ),
	.cordic_x_res_2c_11(\cordinv|cordic_x_res_2c[11]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cord_2c cordinv(
	.cordic_x_res_2c_0(\cordinv|cordic_x_res_2c[0]~q ),
	.cordic_y_res_2c_0(\cordinv|cordic_y_res_2c[0]~q ),
	.cordic_y_res_d_1(\cordinv|cordic_y_res_d[1]~q ),
	.cordic_x_res_d_1(\cordinv|cordic_x_res_d[1]~q ),
	.cordic_y_res_2c_1(\cordinv|cordic_y_res_2c[1]~q ),
	.cordic_x_res_2c_1(\cordinv|cordic_x_res_2c[1]~q ),
	.cordic_y_res_d_2(\cordinv|cordic_y_res_d[2]~q ),
	.cordic_x_res_d_2(\cordinv|cordic_x_res_d[2]~q ),
	.cordic_y_res_2c_2(\cordinv|cordic_y_res_2c[2]~q ),
	.cordic_x_res_2c_2(\cordinv|cordic_x_res_2c[2]~q ),
	.cordic_y_res_d_3(\cordinv|cordic_y_res_d[3]~q ),
	.cordic_x_res_d_3(\cordinv|cordic_x_res_d[3]~q ),
	.cordic_y_res_2c_3(\cordinv|cordic_y_res_2c[3]~q ),
	.cordic_x_res_2c_3(\cordinv|cordic_x_res_2c[3]~q ),
	.cordic_y_res_d_4(\cordinv|cordic_y_res_d[4]~q ),
	.cordic_x_res_d_4(\cordinv|cordic_x_res_d[4]~q ),
	.cordic_y_res_2c_4(\cordinv|cordic_y_res_2c[4]~q ),
	.cordic_x_res_2c_4(\cordinv|cordic_x_res_2c[4]~q ),
	.cordic_y_res_d_5(\cordinv|cordic_y_res_d[5]~q ),
	.cordic_x_res_d_5(\cordinv|cordic_x_res_d[5]~q ),
	.cordic_y_res_2c_5(\cordinv|cordic_y_res_2c[5]~q ),
	.cordic_x_res_2c_5(\cordinv|cordic_x_res_2c[5]~q ),
	.cordic_y_res_d_6(\cordinv|cordic_y_res_d[6]~q ),
	.cordic_x_res_d_6(\cordinv|cordic_x_res_d[6]~q ),
	.cordic_y_res_2c_6(\cordinv|cordic_y_res_2c[6]~q ),
	.cordic_x_res_2c_6(\cordinv|cordic_x_res_2c[6]~q ),
	.cordic_y_res_d_7(\cordinv|cordic_y_res_d[7]~q ),
	.cordic_x_res_d_7(\cordinv|cordic_x_res_d[7]~q ),
	.cordic_y_res_2c_7(\cordinv|cordic_y_res_2c[7]~q ),
	.cordic_x_res_2c_7(\cordinv|cordic_x_res_2c[7]~q ),
	.cordic_y_res_d_8(\cordinv|cordic_y_res_d[8]~q ),
	.cordic_x_res_d_8(\cordinv|cordic_x_res_d[8]~q ),
	.cordic_y_res_2c_8(\cordinv|cordic_y_res_2c[8]~q ),
	.cordic_x_res_2c_8(\cordinv|cordic_x_res_2c[8]~q ),
	.cordic_y_res_d_9(\cordinv|cordic_y_res_d[9]~q ),
	.cordic_x_res_d_9(\cordinv|cordic_x_res_d[9]~q ),
	.cordic_y_res_2c_9(\cordinv|cordic_y_res_2c[9]~q ),
	.cordic_x_res_2c_9(\cordinv|cordic_x_res_2c[9]~q ),
	.cordic_y_res_d_10(\cordinv|cordic_y_res_d[10]~q ),
	.cordic_x_res_d_10(\cordinv|cordic_x_res_d[10]~q ),
	.cordic_y_res_2c_10(\cordinv|cordic_y_res_2c[10]~q ),
	.cordic_x_res_2c_10(\cordinv|cordic_x_res_2c[10]~q ),
	.cordic_y_res_d_11(\cordinv|cordic_y_res_d[11]~q ),
	.cordic_x_res_d_11(\cordinv|cordic_x_res_d[11]~q ),
	.cordic_y_res_2c_11(\cordinv|cordic_y_res_2c[11]~q ),
	.cordic_x_res_2c_11(\cordinv|cordic_x_res_2c[11]~q ),
	.dffe1(\u34|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_0(\u35|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u35|u0|auto_generated|pipeline_dffe[1]~q ),
	.dffe2(\u34|u0|auto_generated|dffe2~q ),
	.pipeline_dffe_2(\u35|u0|auto_generated|pipeline_dffe[2]~q ),
	.dffe3(\u34|u0|auto_generated|dffe3~q ),
	.pipeline_dffe_3(\u35|u0|auto_generated|pipeline_dffe[3]~q ),
	.dffe4(\u34|u0|auto_generated|dffe4~q ),
	.pipeline_dffe_4(\u35|u0|auto_generated|pipeline_dffe[4]~q ),
	.dffe5(\u34|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_5(\u35|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe6(\u34|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_6(\u35|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe7(\u34|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_7(\u35|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe8(\u34|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_8(\u35|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe9(\u34|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_9(\u35|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe10(\u34|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_10(\u35|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe11(\u34|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_11(\u35|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe12(\u34|u0|auto_generated|dffe12~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm_8 u35(
	.pipeline_dffe_0(\u35|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u35|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u35|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u35|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u35|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u35|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u35|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u35|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u35|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u35|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u35|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\u35|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe16(\u33|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_111(\u32|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe12(\u31|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_01(\u32|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_12(\u32|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u32|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u32|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u32|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u32|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u32|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u32|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u32|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u32|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\u32|u0|auto_generated|pipeline_dffe[10]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm_8 u34(
	.dffe1(\u34|u0|auto_generated|dffe1~q ),
	.dffe2(\u34|u0|auto_generated|dffe2~q ),
	.dffe3(\u34|u0|auto_generated|dffe3~q ),
	.dffe4(\u34|u0|auto_generated|dffe4~q ),
	.dffe5(\u34|u0|auto_generated|dffe5~q ),
	.dffe6(\u34|u0|auto_generated|dffe6~q ),
	.dffe7(\u34|u0|auto_generated|dffe7~q ),
	.dffe8(\u34|u0|auto_generated|dffe8~q ),
	.dffe9(\u34|u0|auto_generated|dffe9~q ),
	.dffe10(\u34|u0|auto_generated|dffe10~q ),
	.dffe11(\u34|u0|auto_generated|dffe11~q ),
	.dffe12(\u34|u0|auto_generated|dffe12~q ),
	.dffe16(\u33|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_11(\u32|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe121(\u31|u0|auto_generated|dffe12~q ),
	.dffe13(\u31|u0|auto_generated|dffe1~q ),
	.dffe21(\u31|u0|auto_generated|dffe2~q ),
	.dffe31(\u31|u0|auto_generated|dffe3~q ),
	.dffe41(\u31|u0|auto_generated|dffe4~q ),
	.dffe51(\u31|u0|auto_generated|dffe5~q ),
	.dffe61(\u31|u0|auto_generated|dffe6~q ),
	.dffe71(\u31|u0|auto_generated|dffe7~q ),
	.dffe81(\u31|u0|auto_generated|dffe8~q ),
	.dffe91(\u31|u0|auto_generated|dffe9~q ),
	.dffe101(\u31|u0|auto_generated|dffe10~q ),
	.dffe111(\u31|u0|auto_generated|dffe11~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_zxor_1p_lpm_8 u33(
	.dffe16(\u33|u0|auto_generated|dffe16~q ),
	.dffe161(\u30|u0|auto_generated|dffe16~q ),
	.dffe15(\u30|u0|auto_generated|dffe15~q ),
	.dffe14(\u30|u0|auto_generated|dffe14~q ),
	.dffe13(\u30|u0|auto_generated|dffe13~q ),
	.dffe12(\u30|u0|auto_generated|dffe12~q ),
	.dffe11(\u30|u0|auto_generated|dffe11~q ),
	.dffe10(\u30|u0|auto_generated|dffe10~q ),
	.dffe9(\u30|u0|auto_generated|dffe9~q ),
	.dffe8(\u30|u0|auto_generated|dffe8~q ),
	.dffe7(\u30|u0|auto_generated|dffe7~q ),
	.dffe6(\u30|u0|auto_generated|dffe6~q ),
	.dffe5(\u30|u0|auto_generated|dffe5~q ),
	.dffe4(\u30|u0|auto_generated|dffe4~q ),
	.dffe3(\u30|u0|auto_generated|dffe3~q ),
	.dffe2(\u30|u0|auto_generated|dffe2~q ),
	.dffe1(\u30|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm_7 u32(
	.pipeline_dffe_11(\u32|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_0(\u32|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u32|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u32|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u32|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u32|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u32|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u32|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u32|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u32|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u32|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u32|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe16(\u30|u0|auto_generated|dffe16~q ),
	.dffe12(\u28|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_111(\u29|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_101(\u29|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe11(\u28|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_01(\u29|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_12(\u29|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u29|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u29|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u29|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u29|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u29|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u29|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u29|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u29|u0|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm_7 u31(
	.dffe12(\u31|u0|auto_generated|dffe12~q ),
	.dffe1(\u31|u0|auto_generated|dffe1~q ),
	.dffe2(\u31|u0|auto_generated|dffe2~q ),
	.dffe3(\u31|u0|auto_generated|dffe3~q ),
	.dffe4(\u31|u0|auto_generated|dffe4~q ),
	.dffe5(\u31|u0|auto_generated|dffe5~q ),
	.dffe6(\u31|u0|auto_generated|dffe6~q ),
	.dffe7(\u31|u0|auto_generated|dffe7~q ),
	.dffe8(\u31|u0|auto_generated|dffe8~q ),
	.dffe9(\u31|u0|auto_generated|dffe9~q ),
	.dffe10(\u31|u0|auto_generated|dffe10~q ),
	.dffe11(\u31|u0|auto_generated|dffe11~q ),
	.dffe16(\u30|u0|auto_generated|dffe16~q ),
	.dffe121(\u28|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_11(\u29|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\u29|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe111(\u28|u0|auto_generated|dffe11~q ),
	.dffe13(\u28|u0|auto_generated|dffe1~q ),
	.dffe21(\u28|u0|auto_generated|dffe2~q ),
	.dffe31(\u28|u0|auto_generated|dffe3~q ),
	.dffe41(\u28|u0|auto_generated|dffe4~q ),
	.dffe51(\u28|u0|auto_generated|dffe5~q ),
	.dffe61(\u28|u0|auto_generated|dffe6~q ),
	.dffe71(\u28|u0|auto_generated|dffe7~q ),
	.dffe81(\u28|u0|auto_generated|dffe8~q ),
	.dffe91(\u28|u0|auto_generated|dffe9~q ),
	.dffe101(\u28|u0|auto_generated|dffe10~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_zxor_1p_lpm_7 u30(
	.dffe16(\u30|u0|auto_generated|dffe16~q ),
	.dffe15(\u30|u0|auto_generated|dffe15~q ),
	.dffe14(\u30|u0|auto_generated|dffe14~q ),
	.dffe161(\u27|u0|auto_generated|dffe16~q ),
	.dffe13(\u30|u0|auto_generated|dffe13~q ),
	.dffe12(\u30|u0|auto_generated|dffe12~q ),
	.dffe151(\u27|u0|auto_generated|dffe15~q ),
	.dffe11(\u30|u0|auto_generated|dffe11~q ),
	.dffe141(\u27|u0|auto_generated|dffe14~q ),
	.dffe10(\u30|u0|auto_generated|dffe10~q ),
	.dffe131(\u27|u0|auto_generated|dffe13~q ),
	.dffe9(\u30|u0|auto_generated|dffe9~q ),
	.dffe121(\u27|u0|auto_generated|dffe12~q ),
	.dffe8(\u30|u0|auto_generated|dffe8~q ),
	.dffe111(\u27|u0|auto_generated|dffe11~q ),
	.dffe7(\u30|u0|auto_generated|dffe7~q ),
	.dffe101(\u27|u0|auto_generated|dffe10~q ),
	.dffe6(\u30|u0|auto_generated|dffe6~q ),
	.dffe91(\u27|u0|auto_generated|dffe9~q ),
	.dffe5(\u30|u0|auto_generated|dffe5~q ),
	.dffe81(\u27|u0|auto_generated|dffe8~q ),
	.dffe4(\u30|u0|auto_generated|dffe4~q ),
	.dffe71(\u27|u0|auto_generated|dffe7~q ),
	.dffe3(\u30|u0|auto_generated|dffe3~q ),
	.dffe61(\u27|u0|auto_generated|dffe6~q ),
	.dffe2(\u30|u0|auto_generated|dffe2~q ),
	.dffe51(\u27|u0|auto_generated|dffe5~q ),
	.dffe1(\u30|u0|auto_generated|dffe1~q ),
	.dffe41(\u27|u0|auto_generated|dffe4~q ),
	.dffe31(\u27|u0|auto_generated|dffe3~q ),
	.dffe21(\u27|u0|auto_generated|dffe2~q ),
	.dffe17(\u27|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm_6 u29(
	.pipeline_dffe_11(\u29|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\u29|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_0(\u29|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u29|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u29|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u29|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u29|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u29|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u29|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u29|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u29|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u29|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe16(\u27|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_111(\u26|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe12(\u25|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_91(\u26|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\u26|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe11(\u25|u0|auto_generated|dffe11~q ),
	.dffe10(\u25|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_01(\u26|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_12(\u26|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u26|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u26|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u26|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u26|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u26|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u26|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u26|u0|auto_generated|pipeline_dffe[8]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm_6 u28(
	.dffe12(\u28|u0|auto_generated|dffe12~q ),
	.dffe11(\u28|u0|auto_generated|dffe11~q ),
	.dffe1(\u28|u0|auto_generated|dffe1~q ),
	.dffe2(\u28|u0|auto_generated|dffe2~q ),
	.dffe3(\u28|u0|auto_generated|dffe3~q ),
	.dffe4(\u28|u0|auto_generated|dffe4~q ),
	.dffe5(\u28|u0|auto_generated|dffe5~q ),
	.dffe6(\u28|u0|auto_generated|dffe6~q ),
	.dffe7(\u28|u0|auto_generated|dffe7~q ),
	.dffe8(\u28|u0|auto_generated|dffe8~q ),
	.dffe9(\u28|u0|auto_generated|dffe9~q ),
	.dffe10(\u28|u0|auto_generated|dffe10~q ),
	.dffe16(\u27|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_11(\u26|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe121(\u25|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_9(\u26|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u26|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe111(\u25|u0|auto_generated|dffe11~q ),
	.dffe101(\u25|u0|auto_generated|dffe10~q ),
	.dffe13(\u25|u0|auto_generated|dffe1~q ),
	.dffe21(\u25|u0|auto_generated|dffe2~q ),
	.dffe31(\u25|u0|auto_generated|dffe3~q ),
	.dffe41(\u25|u0|auto_generated|dffe4~q ),
	.dffe51(\u25|u0|auto_generated|dffe5~q ),
	.dffe61(\u25|u0|auto_generated|dffe6~q ),
	.dffe71(\u25|u0|auto_generated|dffe7~q ),
	.dffe81(\u25|u0|auto_generated|dffe8~q ),
	.dffe91(\u25|u0|auto_generated|dffe9~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_zxor_1p_lpm_5 u27(
	.dffe16(\u27|u0|auto_generated|dffe16~q ),
	.dffe15(\u27|u0|auto_generated|dffe15~q ),
	.dffe14(\u27|u0|auto_generated|dffe14~q ),
	.dffe161(\u24|u0|auto_generated|dffe16~q ),
	.dffe13(\u27|u0|auto_generated|dffe13~q ),
	.dffe12(\u27|u0|auto_generated|dffe12~q ),
	.dffe151(\u24|u0|auto_generated|dffe15~q ),
	.dffe11(\u27|u0|auto_generated|dffe11~q ),
	.dffe141(\u24|u0|auto_generated|dffe14~q ),
	.dffe10(\u27|u0|auto_generated|dffe10~q ),
	.dffe131(\u24|u0|auto_generated|dffe13~q ),
	.dffe9(\u27|u0|auto_generated|dffe9~q ),
	.dffe121(\u24|u0|auto_generated|dffe12~q ),
	.dffe8(\u27|u0|auto_generated|dffe8~q ),
	.dffe111(\u24|u0|auto_generated|dffe11~q ),
	.dffe7(\u27|u0|auto_generated|dffe7~q ),
	.dffe101(\u24|u0|auto_generated|dffe10~q ),
	.dffe6(\u27|u0|auto_generated|dffe6~q ),
	.dffe91(\u24|u0|auto_generated|dffe9~q ),
	.dffe5(\u27|u0|auto_generated|dffe5~q ),
	.dffe81(\u24|u0|auto_generated|dffe8~q ),
	.dffe4(\u27|u0|auto_generated|dffe4~q ),
	.dffe71(\u24|u0|auto_generated|dffe7~q ),
	.dffe3(\u27|u0|auto_generated|dffe3~q ),
	.dffe61(\u24|u0|auto_generated|dffe6~q ),
	.dffe2(\u27|u0|auto_generated|dffe2~q ),
	.dffe51(\u24|u0|auto_generated|dffe5~q ),
	.dffe1(\u27|u0|auto_generated|dffe1~q ),
	.dffe41(\u24|u0|auto_generated|dffe4~q ),
	.dffe31(\u24|u0|auto_generated|dffe3~q ),
	.dffe21(\u24|u0|auto_generated|dffe2~q ),
	.dffe17(\u24|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm_5 u26(
	.pipeline_dffe_11(\u26|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_9(\u26|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u26|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe16(\u24|u0|auto_generated|dffe16~q ),
	.dffe12(\u22|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_111(\u23|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_0(\u26|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u26|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u26|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u26|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u26|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u26|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u26|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u26|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u26|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_101(\u23|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe11(\u22|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_81(\u23|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u23|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe10(\u22|u0|auto_generated|dffe10~q ),
	.dffe9(\u22|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_01(\u23|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_12(\u23|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u23|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u23|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u23|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u23|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u23|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u23|u0|auto_generated|pipeline_dffe[7]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm_5 u25(
	.dffe12(\u25|u0|auto_generated|dffe12~q ),
	.dffe11(\u25|u0|auto_generated|dffe11~q ),
	.dffe10(\u25|u0|auto_generated|dffe10~q ),
	.dffe1(\u25|u0|auto_generated|dffe1~q ),
	.dffe16(\u24|u0|auto_generated|dffe16~q ),
	.dffe121(\u22|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_11(\u23|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe2(\u25|u0|auto_generated|dffe2~q ),
	.dffe3(\u25|u0|auto_generated|dffe3~q ),
	.dffe4(\u25|u0|auto_generated|dffe4~q ),
	.dffe5(\u25|u0|auto_generated|dffe5~q ),
	.dffe6(\u25|u0|auto_generated|dffe6~q ),
	.dffe7(\u25|u0|auto_generated|dffe7~q ),
	.dffe8(\u25|u0|auto_generated|dffe8~q ),
	.dffe9(\u25|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_10(\u23|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe111(\u22|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_8(\u23|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u23|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe101(\u22|u0|auto_generated|dffe10~q ),
	.dffe91(\u22|u0|auto_generated|dffe9~q ),
	.dffe13(\u22|u0|auto_generated|dffe1~q ),
	.dffe21(\u22|u0|auto_generated|dffe2~q ),
	.dffe31(\u22|u0|auto_generated|dffe3~q ),
	.dffe41(\u22|u0|auto_generated|dffe4~q ),
	.dffe51(\u22|u0|auto_generated|dffe5~q ),
	.dffe61(\u22|u0|auto_generated|dffe6~q ),
	.dffe71(\u22|u0|auto_generated|dffe7~q ),
	.dffe81(\u22|u0|auto_generated|dffe8~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_zxor_1p_lpm_4 u24(
	.dffe16(\u24|u0|auto_generated|dffe16~q ),
	.dffe15(\u24|u0|auto_generated|dffe15~q ),
	.dffe14(\u24|u0|auto_generated|dffe14~q ),
	.dffe161(\u21|u0|auto_generated|dffe16~q ),
	.dffe13(\u24|u0|auto_generated|dffe13~q ),
	.dffe12(\u24|u0|auto_generated|dffe12~q ),
	.dffe151(\u21|u0|auto_generated|dffe15~q ),
	.dffe11(\u24|u0|auto_generated|dffe11~q ),
	.dffe141(\u21|u0|auto_generated|dffe14~q ),
	.dffe10(\u24|u0|auto_generated|dffe10~q ),
	.dffe131(\u21|u0|auto_generated|dffe13~q ),
	.dffe9(\u24|u0|auto_generated|dffe9~q ),
	.dffe121(\u21|u0|auto_generated|dffe12~q ),
	.dffe8(\u24|u0|auto_generated|dffe8~q ),
	.dffe111(\u21|u0|auto_generated|dffe11~q ),
	.dffe7(\u24|u0|auto_generated|dffe7~q ),
	.dffe101(\u21|u0|auto_generated|dffe10~q ),
	.dffe6(\u24|u0|auto_generated|dffe6~q ),
	.dffe91(\u21|u0|auto_generated|dffe9~q ),
	.dffe5(\u24|u0|auto_generated|dffe5~q ),
	.dffe81(\u21|u0|auto_generated|dffe8~q ),
	.dffe4(\u24|u0|auto_generated|dffe4~q ),
	.dffe71(\u21|u0|auto_generated|dffe7~q ),
	.dffe3(\u24|u0|auto_generated|dffe3~q ),
	.dffe61(\u21|u0|auto_generated|dffe6~q ),
	.dffe2(\u24|u0|auto_generated|dffe2~q ),
	.dffe51(\u21|u0|auto_generated|dffe5~q ),
	.dffe1(\u24|u0|auto_generated|dffe1~q ),
	.dffe41(\u21|u0|auto_generated|dffe4~q ),
	.dffe31(\u21|u0|auto_generated|dffe3~q ),
	.dffe21(\u21|u0|auto_generated|dffe2~q ),
	.dffe17(\u21|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm_4 u23(
	.pipeline_dffe_11(\u23|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\u23|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_8(\u23|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u23|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe16(\u21|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_111(\u20|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe12(\u19|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_0(\u23|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u23|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u23|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u23|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u23|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u23|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u23|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u23|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe11(\u19|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_101(\u20|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe10(\u19|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_91(\u20|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_71(\u20|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u20|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe9(\u19|u0|auto_generated|dffe9~q ),
	.dffe8(\u19|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_01(\u20|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_12(\u20|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u20|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u20|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u20|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u20|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u20|u0|auto_generated|pipeline_dffe[6]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm_4 u22(
	.dffe12(\u22|u0|auto_generated|dffe12~q ),
	.dffe11(\u22|u0|auto_generated|dffe11~q ),
	.dffe16(\u21|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_11(\u20|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe10(\u22|u0|auto_generated|dffe10~q ),
	.dffe121(\u19|u0|auto_generated|dffe12~q ),
	.dffe9(\u22|u0|auto_generated|dffe9~q ),
	.dffe1(\u22|u0|auto_generated|dffe1~q ),
	.dffe2(\u22|u0|auto_generated|dffe2~q ),
	.dffe3(\u22|u0|auto_generated|dffe3~q ),
	.dffe4(\u22|u0|auto_generated|dffe4~q ),
	.dffe5(\u22|u0|auto_generated|dffe5~q ),
	.dffe6(\u22|u0|auto_generated|dffe6~q ),
	.dffe7(\u22|u0|auto_generated|dffe7~q ),
	.dffe8(\u22|u0|auto_generated|dffe8~q ),
	.dffe111(\u19|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_10(\u20|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe101(\u19|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_9(\u20|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_7(\u20|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u20|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe91(\u19|u0|auto_generated|dffe9~q ),
	.dffe81(\u19|u0|auto_generated|dffe8~q ),
	.dffe13(\u19|u0|auto_generated|dffe1~q ),
	.dffe21(\u19|u0|auto_generated|dffe2~q ),
	.dffe31(\u19|u0|auto_generated|dffe3~q ),
	.dffe41(\u19|u0|auto_generated|dffe4~q ),
	.dffe51(\u19|u0|auto_generated|dffe5~q ),
	.dffe61(\u19|u0|auto_generated|dffe6~q ),
	.dffe71(\u19|u0|auto_generated|dffe7~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_zxor_1p_lpm_3 u21(
	.dffe16(\u21|u0|auto_generated|dffe16~q ),
	.dffe15(\u21|u0|auto_generated|dffe15~q ),
	.dffe14(\u21|u0|auto_generated|dffe14~q ),
	.dffe161(\u18|u0|auto_generated|dffe16~q ),
	.dffe13(\u21|u0|auto_generated|dffe13~q ),
	.dffe12(\u21|u0|auto_generated|dffe12~q ),
	.dffe151(\u18|u0|auto_generated|dffe15~q ),
	.dffe11(\u21|u0|auto_generated|dffe11~q ),
	.dffe141(\u18|u0|auto_generated|dffe14~q ),
	.dffe10(\u21|u0|auto_generated|dffe10~q ),
	.dffe131(\u18|u0|auto_generated|dffe13~q ),
	.dffe9(\u21|u0|auto_generated|dffe9~q ),
	.dffe121(\u18|u0|auto_generated|dffe12~q ),
	.dffe8(\u21|u0|auto_generated|dffe8~q ),
	.dffe111(\u18|u0|auto_generated|dffe11~q ),
	.dffe7(\u21|u0|auto_generated|dffe7~q ),
	.dffe101(\u18|u0|auto_generated|dffe10~q ),
	.dffe6(\u21|u0|auto_generated|dffe6~q ),
	.dffe91(\u18|u0|auto_generated|dffe9~q ),
	.dffe5(\u21|u0|auto_generated|dffe5~q ),
	.dffe81(\u18|u0|auto_generated|dffe8~q ),
	.dffe4(\u21|u0|auto_generated|dffe4~q ),
	.dffe71(\u18|u0|auto_generated|dffe7~q ),
	.dffe3(\u21|u0|auto_generated|dffe3~q ),
	.dffe61(\u18|u0|auto_generated|dffe6~q ),
	.dffe2(\u21|u0|auto_generated|dffe2~q ),
	.dffe51(\u18|u0|auto_generated|dffe5~q ),
	.dffe1(\u21|u0|auto_generated|dffe1~q ),
	.dffe41(\u18|u0|auto_generated|dffe4~q ),
	.dffe31(\u18|u0|auto_generated|dffe3~q ),
	.dffe21(\u18|u0|auto_generated|dffe2~q ),
	.dffe17(\u18|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm_3 u20(
	.pipeline_dffe_11(\u20|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\u20|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe16(\u18|u0|auto_generated|dffe16~q ),
	.dffe12(\u16|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_9(\u20|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_111(\u17|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_7(\u20|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u20|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_101(\u17|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe11(\u16|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_0(\u20|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u20|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u20|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u20|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u20|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u20|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u20|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_91(\u17|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe10(\u16|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_81(\u17|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe9(\u16|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_61(\u17|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u17|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe8(\u16|u0|auto_generated|dffe8~q ),
	.dffe7(\u16|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_01(\u17|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_12(\u17|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u17|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u17|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u17|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u17|u0|auto_generated|pipeline_dffe[5]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm_3 u19(
	.dffe12(\u19|u0|auto_generated|dffe12~q ),
	.dffe11(\u19|u0|auto_generated|dffe11~q ),
	.dffe16(\u18|u0|auto_generated|dffe16~q ),
	.dffe10(\u19|u0|auto_generated|dffe10~q ),
	.dffe121(\u16|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_11(\u17|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe9(\u19|u0|auto_generated|dffe9~q ),
	.dffe8(\u19|u0|auto_generated|dffe8~q ),
	.dffe1(\u19|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_10(\u17|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe111(\u16|u0|auto_generated|dffe11~q ),
	.dffe2(\u19|u0|auto_generated|dffe2~q ),
	.dffe3(\u19|u0|auto_generated|dffe3~q ),
	.dffe4(\u19|u0|auto_generated|dffe4~q ),
	.dffe5(\u19|u0|auto_generated|dffe5~q ),
	.dffe6(\u19|u0|auto_generated|dffe6~q ),
	.dffe7(\u19|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_9(\u17|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe101(\u16|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_8(\u17|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe91(\u16|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_6(\u17|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u17|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe81(\u16|u0|auto_generated|dffe8~q ),
	.dffe71(\u16|u0|auto_generated|dffe7~q ),
	.dffe13(\u16|u0|auto_generated|dffe1~q ),
	.dffe21(\u16|u0|auto_generated|dffe2~q ),
	.dffe31(\u16|u0|auto_generated|dffe3~q ),
	.dffe41(\u16|u0|auto_generated|dffe4~q ),
	.dffe51(\u16|u0|auto_generated|dffe5~q ),
	.dffe61(\u16|u0|auto_generated|dffe6~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_zxor_1p_lpm_2 u18(
	.dffe16(\u18|u0|auto_generated|dffe16~q ),
	.dffe15(\u18|u0|auto_generated|dffe15~q ),
	.dffe14(\u18|u0|auto_generated|dffe14~q ),
	.dffe161(\u15|u0|auto_generated|dffe16~q ),
	.dffe13(\u18|u0|auto_generated|dffe13~q ),
	.dffe12(\u18|u0|auto_generated|dffe12~q ),
	.dffe151(\u15|u0|auto_generated|dffe15~q ),
	.dffe11(\u18|u0|auto_generated|dffe11~q ),
	.dffe141(\u15|u0|auto_generated|dffe14~q ),
	.dffe10(\u18|u0|auto_generated|dffe10~q ),
	.dffe131(\u15|u0|auto_generated|dffe13~q ),
	.dffe9(\u18|u0|auto_generated|dffe9~q ),
	.dffe121(\u15|u0|auto_generated|dffe12~q ),
	.dffe8(\u18|u0|auto_generated|dffe8~q ),
	.dffe111(\u15|u0|auto_generated|dffe11~q ),
	.dffe7(\u18|u0|auto_generated|dffe7~q ),
	.dffe101(\u15|u0|auto_generated|dffe10~q ),
	.dffe6(\u18|u0|auto_generated|dffe6~q ),
	.dffe91(\u15|u0|auto_generated|dffe9~q ),
	.dffe5(\u18|u0|auto_generated|dffe5~q ),
	.dffe81(\u15|u0|auto_generated|dffe8~q ),
	.dffe4(\u18|u0|auto_generated|dffe4~q ),
	.dffe71(\u15|u0|auto_generated|dffe7~q ),
	.dffe3(\u18|u0|auto_generated|dffe3~q ),
	.dffe61(\u15|u0|auto_generated|dffe6~q ),
	.dffe2(\u18|u0|auto_generated|dffe2~q ),
	.dffe51(\u15|u0|auto_generated|dffe5~q ),
	.dffe1(\u18|u0|auto_generated|dffe1~q ),
	.dffe41(\u15|u0|auto_generated|dffe4~q ),
	.dffe31(\u15|u0|auto_generated|dffe3~q ),
	.dffe21(\u15|u0|auto_generated|dffe2~q ),
	.dffe17(\u15|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm_2 u17(
	.pipeline_dffe_11(\u17|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\u17|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe16(\u15|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_9(\u17|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_111(\u14|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe12(\u13|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_8(\u17|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_6(\u17|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u17|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe11(\u13|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_101(\u14|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe10(\u13|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_91(\u14|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_0(\u17|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u17|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u17|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u17|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u17|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u17|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe9(\u13|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_81(\u14|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe8(\u13|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_71(\u14|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_51(\u14|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u14|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe7(\u13|u0|auto_generated|dffe7~q ),
	.dffe6(\u13|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_01(\u14|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_12(\u14|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u14|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u14|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u14|u0|auto_generated|pipeline_dffe[4]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm_2 u16(
	.dffe12(\u16|u0|auto_generated|dffe12~q ),
	.dffe11(\u16|u0|auto_generated|dffe11~q ),
	.dffe16(\u15|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_11(\u14|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe10(\u16|u0|auto_generated|dffe10~q ),
	.dffe121(\u13|u0|auto_generated|dffe12~q ),
	.dffe9(\u16|u0|auto_generated|dffe9~q ),
	.dffe111(\u13|u0|auto_generated|dffe11~q ),
	.dffe8(\u16|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_10(\u14|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe7(\u16|u0|auto_generated|dffe7~q ),
	.dffe1(\u16|u0|auto_generated|dffe1~q ),
	.dffe101(\u13|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_9(\u14|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe2(\u16|u0|auto_generated|dffe2~q ),
	.dffe3(\u16|u0|auto_generated|dffe3~q ),
	.dffe4(\u16|u0|auto_generated|dffe4~q ),
	.dffe5(\u16|u0|auto_generated|dffe5~q ),
	.dffe6(\u16|u0|auto_generated|dffe6~q ),
	.dffe91(\u13|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_8(\u14|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe81(\u13|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_7(\u14|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_5(\u14|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u14|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe71(\u13|u0|auto_generated|dffe7~q ),
	.dffe61(\u13|u0|auto_generated|dffe6~q ),
	.dffe13(\u13|u0|auto_generated|dffe1~q ),
	.dffe21(\u13|u0|auto_generated|dffe2~q ),
	.dffe31(\u13|u0|auto_generated|dffe3~q ),
	.dffe41(\u13|u0|auto_generated|dffe4~q ),
	.dffe51(\u13|u0|auto_generated|dffe5~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_zxor_1p_lpm_1 u15(
	.dffe16(\u15|u0|auto_generated|dffe16~q ),
	.dffe15(\u15|u0|auto_generated|dffe15~q ),
	.dffe14(\u15|u0|auto_generated|dffe14~q ),
	.dffe161(\u12|u0|auto_generated|dffe16~q ),
	.dffe13(\u15|u0|auto_generated|dffe13~q ),
	.dffe12(\u15|u0|auto_generated|dffe12~q ),
	.dffe151(\u12|u0|auto_generated|dffe15~q ),
	.dffe11(\u15|u0|auto_generated|dffe11~q ),
	.dffe141(\u12|u0|auto_generated|dffe14~q ),
	.dffe10(\u15|u0|auto_generated|dffe10~q ),
	.dffe131(\u12|u0|auto_generated|dffe13~q ),
	.dffe9(\u15|u0|auto_generated|dffe9~q ),
	.dffe121(\u12|u0|auto_generated|dffe12~q ),
	.dffe8(\u15|u0|auto_generated|dffe8~q ),
	.dffe111(\u12|u0|auto_generated|dffe11~q ),
	.dffe7(\u15|u0|auto_generated|dffe7~q ),
	.dffe101(\u12|u0|auto_generated|dffe10~q ),
	.dffe6(\u15|u0|auto_generated|dffe6~q ),
	.dffe91(\u12|u0|auto_generated|dffe9~q ),
	.dffe5(\u15|u0|auto_generated|dffe5~q ),
	.dffe81(\u12|u0|auto_generated|dffe8~q ),
	.dffe4(\u15|u0|auto_generated|dffe4~q ),
	.dffe71(\u12|u0|auto_generated|dffe7~q ),
	.dffe3(\u15|u0|auto_generated|dffe3~q ),
	.dffe61(\u12|u0|auto_generated|dffe6~q ),
	.dffe2(\u15|u0|auto_generated|dffe2~q ),
	.dffe51(\u12|u0|auto_generated|dffe5~q ),
	.dffe1(\u15|u0|auto_generated|dffe1~q ),
	.dffe41(\u12|u0|auto_generated|dffe4~q ),
	.dffe31(\u12|u0|auto_generated|dffe3~q ),
	.dffe21(\u12|u0|auto_generated|dffe2~q ),
	.dffe17(\u12|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm_1 u14(
	.pipeline_dffe_11(\u14|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\u14|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe16(\u12|u0|auto_generated|dffe16~q ),
	.dffe12(\u10|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_9(\u14|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_111(\u11|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_8(\u14|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_101(\u11|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_7(\u14|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe11(\u10|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_5(\u14|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u14|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_91(\u11|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe10(\u10|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_81(\u11|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe9(\u10|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_0(\u14|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u14|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u14|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u14|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u14|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_71(\u11|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe8(\u10|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_61(\u11|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe7(\u10|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_41(\u11|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u11|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe6(\u10|u0|auto_generated|dffe6~q ),
	.dffe5(\u10|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_01(\u11|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_12(\u11|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u11|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u11|u0|auto_generated|pipeline_dffe[3]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm_1 u13(
	.dffe12(\u13|u0|auto_generated|dffe12~q ),
	.dffe11(\u13|u0|auto_generated|dffe11~q ),
	.dffe16(\u12|u0|auto_generated|dffe16~q ),
	.dffe10(\u13|u0|auto_generated|dffe10~q ),
	.dffe121(\u10|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_11(\u11|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe9(\u13|u0|auto_generated|dffe9~q ),
	.dffe8(\u13|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_10(\u11|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe111(\u10|u0|auto_generated|dffe11~q ),
	.dffe7(\u13|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_9(\u11|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe101(\u10|u0|auto_generated|dffe10~q ),
	.dffe6(\u13|u0|auto_generated|dffe6~q ),
	.dffe1(\u13|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_8(\u11|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe91(\u10|u0|auto_generated|dffe9~q ),
	.dffe2(\u13|u0|auto_generated|dffe2~q ),
	.dffe3(\u13|u0|auto_generated|dffe3~q ),
	.dffe4(\u13|u0|auto_generated|dffe4~q ),
	.dffe5(\u13|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_7(\u11|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe81(\u10|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_6(\u11|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe71(\u10|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_4(\u11|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u11|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe61(\u10|u0|auto_generated|dffe6~q ),
	.dffe51(\u10|u0|auto_generated|dffe5~q ),
	.dffe13(\u10|u0|auto_generated|dffe1~q ),
	.dffe21(\u10|u0|auto_generated|dffe2~q ),
	.dffe31(\u10|u0|auto_generated|dffe3~q ),
	.dffe41(\u10|u0|auto_generated|dffe4~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_zxor_1p_lpm u12(
	.dffe16(\u12|u0|auto_generated|dffe16~q ),
	.dffe15(\u12|u0|auto_generated|dffe15~q ),
	.dffe14(\u12|u0|auto_generated|dffe14~q ),
	.dffe161(\u9|u0|auto_generated|dffe16~q ),
	.dffe13(\u12|u0|auto_generated|dffe13~q ),
	.dffe12(\u12|u0|auto_generated|dffe12~q ),
	.dffe151(\u9|u0|auto_generated|dffe15~q ),
	.dffe11(\u12|u0|auto_generated|dffe11~q ),
	.dffe141(\u9|u0|auto_generated|dffe14~q ),
	.dffe10(\u12|u0|auto_generated|dffe10~q ),
	.dffe131(\u9|u0|auto_generated|dffe13~q ),
	.dffe9(\u12|u0|auto_generated|dffe9~q ),
	.dffe121(\u9|u0|auto_generated|dffe12~q ),
	.dffe8(\u12|u0|auto_generated|dffe8~q ),
	.dffe111(\u9|u0|auto_generated|dffe11~q ),
	.dffe7(\u12|u0|auto_generated|dffe7~q ),
	.dffe101(\u9|u0|auto_generated|dffe10~q ),
	.dffe6(\u12|u0|auto_generated|dffe6~q ),
	.dffe91(\u9|u0|auto_generated|dffe9~q ),
	.dffe5(\u12|u0|auto_generated|dffe5~q ),
	.dffe81(\u9|u0|auto_generated|dffe8~q ),
	.dffe4(\u12|u0|auto_generated|dffe4~q ),
	.dffe71(\u9|u0|auto_generated|dffe7~q ),
	.dffe3(\u12|u0|auto_generated|dffe3~q ),
	.dffe61(\u9|u0|auto_generated|dffe6~q ),
	.dffe2(\u12|u0|auto_generated|dffe2~q ),
	.dffe51(\u9|u0|auto_generated|dffe5~q ),
	.dffe1(\u12|u0|auto_generated|dffe1~q ),
	.dffe41(\u9|u0|auto_generated|dffe4~q ),
	.dffe31(\u9|u0|auto_generated|dffe3~q ),
	.dffe21(\u9|u0|auto_generated|dffe2~q ),
	.dffe17(\u9|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_axor_1p_lpm u11(
	.pipeline_dffe_11(\u11|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\u11|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe16(\u9|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_9(\u11|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_111(\u8|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe12(\u7|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_8(\u11|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\u11|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe11(\u7|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_101(\u8|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_6(\u11|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe10(\u7|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_91(\u8|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_4(\u11|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u11|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe9(\u7|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_81(\u8|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe8(\u7|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_71(\u8|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_0(\u11|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u11|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u11|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u11|u0|auto_generated|pipeline_dffe[3]~q ),
	.dffe7(\u7|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_61(\u8|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe6(\u7|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_51(\u8|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_31(\u8|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u8|u0|auto_generated|pipeline_dffe[4]~q ),
	.dffe5(\u7|u0|auto_generated|dffe5~q ),
	.dffe4(\u7|u0|auto_generated|dffe4~q ),
	.pipeline_dffe_01(\u8|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_12(\u8|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u8|u0|auto_generated|pipeline_dffe[2]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_cordic_sxor_1p_lpm u10(
	.dffe12(\u10|u0|auto_generated|dffe12~q ),
	.dffe11(\u10|u0|auto_generated|dffe11~q ),
	.dffe16(\u9|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_11(\u8|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe10(\u10|u0|auto_generated|dffe10~q ),
	.dffe121(\u7|u0|auto_generated|dffe12~q ),
	.dffe9(\u10|u0|auto_generated|dffe9~q ),
	.dffe111(\u7|u0|auto_generated|dffe11~q ),
	.dffe8(\u10|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_10(\u8|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe101(\u7|u0|auto_generated|dffe10~q ),
	.dffe7(\u10|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_9(\u8|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe91(\u7|u0|auto_generated|dffe9~q ),
	.dffe6(\u10|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_8(\u8|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe5(\u10|u0|auto_generated|dffe5~q ),
	.dffe1(\u10|u0|auto_generated|dffe1~q ),
	.dffe81(\u7|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_7(\u8|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe2(\u10|u0|auto_generated|dffe2~q ),
	.dffe3(\u10|u0|auto_generated|dffe3~q ),
	.dffe4(\u10|u0|auto_generated|dffe4~q ),
	.dffe71(\u7|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_6(\u8|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe61(\u7|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_5(\u8|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_3(\u8|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u8|u0|auto_generated|pipeline_dffe[4]~q ),
	.dffe51(\u7|u0|auto_generated|dffe5~q ),
	.dffe41(\u7|u0|auto_generated|dffe4~q ),
	.dffe13(\u7|u0|auto_generated|dffe1~q ),
	.dffe21(\u7|u0|auto_generated|dffe2~q ),
	.dffe31(\u7|u0|auto_generated|dffe3~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

NCO_Lab3_asj_nco_isdr ux710isdr(
	.data_ready1(data_ready),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_asj_altqmcpipe (
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_20,
	pipeline_dffe_19,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	clk,
	reset_n,
	clken,
	phi_inc_i_30,
	phi_inc_i_31,
	phi_inc_i_29,
	phi_inc_i_28,
	phi_inc_i_27,
	phi_inc_i_26,
	phi_inc_i_25,
	phi_inc_i_24,
	phi_inc_i_23,
	phi_inc_i_22,
	phi_inc_i_21,
	phi_inc_i_20,
	phi_inc_i_19,
	phi_inc_i_18,
	phi_inc_i_17,
	phi_inc_i_16,
	phi_inc_i_15,
	phi_inc_i_14,
	phi_inc_i_13,
	phi_inc_i_12,
	phi_inc_i_11,
	phi_inc_i_10,
	phi_inc_i_9,
	phi_inc_i_8,
	phi_inc_i_7,
	phi_inc_i_6,
	phi_inc_i_5,
	phi_inc_i_4,
	phi_inc_i_3,
	phi_inc_i_2,
	phi_inc_i_1,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
output 	pipeline_dffe_29;
output 	pipeline_dffe_28;
output 	pipeline_dffe_27;
output 	pipeline_dffe_26;
output 	pipeline_dffe_25;
output 	pipeline_dffe_24;
output 	pipeline_dffe_23;
output 	pipeline_dffe_22;
output 	pipeline_dffe_21;
output 	pipeline_dffe_20;
output 	pipeline_dffe_19;
output 	pipeline_dffe_18;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
input 	clk;
input 	reset_n;
input 	clken;
input 	phi_inc_i_30;
input 	phi_inc_i_31;
input 	phi_inc_i_29;
input 	phi_inc_i_28;
input 	phi_inc_i_27;
input 	phi_inc_i_26;
input 	phi_inc_i_25;
input 	phi_inc_i_24;
input 	phi_inc_i_23;
input 	phi_inc_i_22;
input 	phi_inc_i_21;
input 	phi_inc_i_20;
input 	phi_inc_i_19;
input 	phi_inc_i_18;
input 	phi_inc_i_17;
input 	phi_inc_i_16;
input 	phi_inc_i_15;
input 	phi_inc_i_14;
input 	phi_inc_i_13;
input 	phi_inc_i_12;
input 	phi_inc_i_11;
input 	phi_inc_i_10;
input 	phi_inc_i_9;
input 	phi_inc_i_8;
input 	phi_inc_i_7;
input 	phi_inc_i_6;
input 	phi_inc_i_5;
input 	phi_inc_i_4;
input 	phi_inc_i_3;
input 	phi_inc_i_2;
input 	phi_inc_i_1;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \phi_int_arr_reg[30]~q ;
wire \phi_int_arr_reg[31]~q ;
wire \phi_int_arr_reg[29]~q ;
wire \phi_int_arr_reg[28]~q ;
wire \phi_int_arr_reg[27]~q ;
wire \phi_int_arr_reg[26]~q ;
wire \phi_int_arr_reg[25]~q ;
wire \phi_int_arr_reg[24]~q ;
wire \phi_int_arr_reg[23]~q ;
wire \phi_int_arr_reg[22]~q ;
wire \phi_int_arr_reg[21]~q ;
wire \phi_int_arr_reg[20]~q ;
wire \phi_int_arr_reg[19]~q ;
wire \phi_int_arr_reg[18]~q ;
wire \phi_int_arr_reg[17]~q ;
wire \phi_int_arr_reg[16]~q ;
wire \phi_int_arr_reg[15]~q ;
wire \phi_int_arr_reg[14]~q ;
wire \phi_int_arr_reg[13]~q ;
wire \phi_int_arr_reg[12]~q ;
wire \phi_int_arr_reg[11]~q ;
wire \phi_int_arr_reg[10]~q ;
wire \phi_int_arr_reg[9]~q ;
wire \phi_int_arr_reg[8]~q ;
wire \phi_int_arr_reg[7]~q ;
wire \phi_int_arr_reg[6]~q ;
wire \phi_int_arr_reg[5]~q ;
wire \phi_int_arr_reg[4]~q ;
wire \phi_int_arr_reg[3]~q ;
wire \phi_int_arr_reg[2]~q ;
wire \phi_int_arr_reg[1]~q ;
wire \phi_int_arr_reg[0]~q ;


NCO_Lab3_lpm_add_sub_1 acc(
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_29(pipeline_dffe_29),
	.phi_int_arr_reg_30(\phi_int_arr_reg[30]~q ),
	.pipeline_dffe_28(pipeline_dffe_28),
	.phi_int_arr_reg_31(\phi_int_arr_reg[31]~q ),
	.phi_int_arr_reg_29(\phi_int_arr_reg[29]~q ),
	.pipeline_dffe_27(pipeline_dffe_27),
	.phi_int_arr_reg_28(\phi_int_arr_reg[28]~q ),
	.pipeline_dffe_26(pipeline_dffe_26),
	.phi_int_arr_reg_27(\phi_int_arr_reg[27]~q ),
	.pipeline_dffe_25(pipeline_dffe_25),
	.phi_int_arr_reg_26(\phi_int_arr_reg[26]~q ),
	.pipeline_dffe_24(pipeline_dffe_24),
	.phi_int_arr_reg_25(\phi_int_arr_reg[25]~q ),
	.pipeline_dffe_23(pipeline_dffe_23),
	.phi_int_arr_reg_24(\phi_int_arr_reg[24]~q ),
	.pipeline_dffe_22(pipeline_dffe_22),
	.phi_int_arr_reg_23(\phi_int_arr_reg[23]~q ),
	.pipeline_dffe_21(pipeline_dffe_21),
	.phi_int_arr_reg_22(\phi_int_arr_reg[22]~q ),
	.pipeline_dffe_20(pipeline_dffe_20),
	.phi_int_arr_reg_21(\phi_int_arr_reg[21]~q ),
	.pipeline_dffe_19(pipeline_dffe_19),
	.phi_int_arr_reg_20(\phi_int_arr_reg[20]~q ),
	.pipeline_dffe_18(pipeline_dffe_18),
	.phi_int_arr_reg_19(\phi_int_arr_reg[19]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.phi_int_arr_reg_18(\phi_int_arr_reg[18]~q ),
	.pipeline_dffe_16(pipeline_dffe_16),
	.phi_int_arr_reg_17(\phi_int_arr_reg[17]~q ),
	.pipeline_dffe_15(pipeline_dffe_15),
	.phi_int_arr_reg_16(\phi_int_arr_reg[16]~q ),
	.pipeline_dffe_14(pipeline_dffe_14),
	.phi_int_arr_reg_15(\phi_int_arr_reg[15]~q ),
	.pipeline_dffe_13(pipeline_dffe_13),
	.phi_int_arr_reg_14(\phi_int_arr_reg[14]~q ),
	.pipeline_dffe_12(pipeline_dffe_12),
	.phi_int_arr_reg_13(\phi_int_arr_reg[13]~q ),
	.pipeline_dffe_11(pipeline_dffe_11),
	.phi_int_arr_reg_12(\phi_int_arr_reg[12]~q ),
	.phi_int_arr_reg_11(\phi_int_arr_reg[11]~q ),
	.phi_int_arr_reg_10(\phi_int_arr_reg[10]~q ),
	.phi_int_arr_reg_9(\phi_int_arr_reg[9]~q ),
	.phi_int_arr_reg_8(\phi_int_arr_reg[8]~q ),
	.phi_int_arr_reg_7(\phi_int_arr_reg[7]~q ),
	.phi_int_arr_reg_6(\phi_int_arr_reg[6]~q ),
	.phi_int_arr_reg_5(\phi_int_arr_reg[5]~q ),
	.phi_int_arr_reg_4(\phi_int_arr_reg[4]~q ),
	.phi_int_arr_reg_3(\phi_int_arr_reg[3]~q ),
	.phi_int_arr_reg_2(\phi_int_arr_reg[2]~q ),
	.phi_int_arr_reg_1(\phi_int_arr_reg[1]~q ),
	.phi_int_arr_reg_0(\phi_int_arr_reg[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \phi_int_arr_reg[30] (
	.clk(clk),
	.d(phi_inc_i_30),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[30]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[30] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[30] .power_up = "low";

dffeas \phi_int_arr_reg[31] (
	.clk(clk),
	.d(phi_inc_i_31),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[31]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[31] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[31] .power_up = "low";

dffeas \phi_int_arr_reg[29] (
	.clk(clk),
	.d(phi_inc_i_29),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[29]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[29] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[29] .power_up = "low";

dffeas \phi_int_arr_reg[28] (
	.clk(clk),
	.d(phi_inc_i_28),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[28]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[28] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[28] .power_up = "low";

dffeas \phi_int_arr_reg[27] (
	.clk(clk),
	.d(phi_inc_i_27),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[27]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[27] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[27] .power_up = "low";

dffeas \phi_int_arr_reg[26] (
	.clk(clk),
	.d(phi_inc_i_26),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[26]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[26] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[26] .power_up = "low";

dffeas \phi_int_arr_reg[25] (
	.clk(clk),
	.d(phi_inc_i_25),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[25]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[25] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[25] .power_up = "low";

dffeas \phi_int_arr_reg[24] (
	.clk(clk),
	.d(phi_inc_i_24),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[24]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[24] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[24] .power_up = "low";

dffeas \phi_int_arr_reg[23] (
	.clk(clk),
	.d(phi_inc_i_23),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[23]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[23] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[23] .power_up = "low";

dffeas \phi_int_arr_reg[22] (
	.clk(clk),
	.d(phi_inc_i_22),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[22]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[22] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[22] .power_up = "low";

dffeas \phi_int_arr_reg[21] (
	.clk(clk),
	.d(phi_inc_i_21),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[21]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[21] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[21] .power_up = "low";

dffeas \phi_int_arr_reg[20] (
	.clk(clk),
	.d(phi_inc_i_20),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[20]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[20] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[20] .power_up = "low";

dffeas \phi_int_arr_reg[19] (
	.clk(clk),
	.d(phi_inc_i_19),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[19]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[19] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[19] .power_up = "low";

dffeas \phi_int_arr_reg[18] (
	.clk(clk),
	.d(phi_inc_i_18),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[18]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[18] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[18] .power_up = "low";

dffeas \phi_int_arr_reg[17] (
	.clk(clk),
	.d(phi_inc_i_17),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[17]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[17] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[17] .power_up = "low";

dffeas \phi_int_arr_reg[16] (
	.clk(clk),
	.d(phi_inc_i_16),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[16]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[16] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[16] .power_up = "low";

dffeas \phi_int_arr_reg[15] (
	.clk(clk),
	.d(phi_inc_i_15),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[15]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[15] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[15] .power_up = "low";

dffeas \phi_int_arr_reg[14] (
	.clk(clk),
	.d(phi_inc_i_14),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[14]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[14] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[14] .power_up = "low";

dffeas \phi_int_arr_reg[13] (
	.clk(clk),
	.d(phi_inc_i_13),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[13]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[13] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[13] .power_up = "low";

dffeas \phi_int_arr_reg[12] (
	.clk(clk),
	.d(phi_inc_i_12),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[12]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[12] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[12] .power_up = "low";

dffeas \phi_int_arr_reg[11] (
	.clk(clk),
	.d(phi_inc_i_11),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[11]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[11] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[11] .power_up = "low";

dffeas \phi_int_arr_reg[10] (
	.clk(clk),
	.d(phi_inc_i_10),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[10]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[10] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[10] .power_up = "low";

dffeas \phi_int_arr_reg[9] (
	.clk(clk),
	.d(phi_inc_i_9),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[9]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[9] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[9] .power_up = "low";

dffeas \phi_int_arr_reg[8] (
	.clk(clk),
	.d(phi_inc_i_8),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[8]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[8] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[8] .power_up = "low";

dffeas \phi_int_arr_reg[7] (
	.clk(clk),
	.d(phi_inc_i_7),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[7]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[7] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[7] .power_up = "low";

dffeas \phi_int_arr_reg[6] (
	.clk(clk),
	.d(phi_inc_i_6),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[6]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[6] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[6] .power_up = "low";

dffeas \phi_int_arr_reg[5] (
	.clk(clk),
	.d(phi_inc_i_5),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[5]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[5] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[5] .power_up = "low";

dffeas \phi_int_arr_reg[4] (
	.clk(clk),
	.d(phi_inc_i_4),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[4]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[4] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[4] .power_up = "low";

dffeas \phi_int_arr_reg[3] (
	.clk(clk),
	.d(phi_inc_i_3),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[3]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[3] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[3] .power_up = "low";

dffeas \phi_int_arr_reg[2] (
	.clk(clk),
	.d(phi_inc_i_2),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[2]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[2] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[2] .power_up = "low";

dffeas \phi_int_arr_reg[1] (
	.clk(clk),
	.d(phi_inc_i_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[1]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[1] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[1] .power_up = "low";

dffeas \phi_int_arr_reg[0] (
	.clk(clk),
	.d(phi_inc_i_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\phi_int_arr_reg[0]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[0] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[0] .power_up = "low";

endmodule

module NCO_Lab3_lpm_add_sub_1 (
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_29,
	phi_int_arr_reg_30,
	pipeline_dffe_28,
	phi_int_arr_reg_31,
	phi_int_arr_reg_29,
	pipeline_dffe_27,
	phi_int_arr_reg_28,
	pipeline_dffe_26,
	phi_int_arr_reg_27,
	pipeline_dffe_25,
	phi_int_arr_reg_26,
	pipeline_dffe_24,
	phi_int_arr_reg_25,
	pipeline_dffe_23,
	phi_int_arr_reg_24,
	pipeline_dffe_22,
	phi_int_arr_reg_23,
	pipeline_dffe_21,
	phi_int_arr_reg_22,
	pipeline_dffe_20,
	phi_int_arr_reg_21,
	pipeline_dffe_19,
	phi_int_arr_reg_20,
	pipeline_dffe_18,
	phi_int_arr_reg_19,
	pipeline_dffe_17,
	phi_int_arr_reg_18,
	pipeline_dffe_16,
	phi_int_arr_reg_17,
	pipeline_dffe_15,
	phi_int_arr_reg_16,
	pipeline_dffe_14,
	phi_int_arr_reg_15,
	pipeline_dffe_13,
	phi_int_arr_reg_14,
	pipeline_dffe_12,
	phi_int_arr_reg_13,
	pipeline_dffe_11,
	phi_int_arr_reg_12,
	phi_int_arr_reg_11,
	phi_int_arr_reg_10,
	phi_int_arr_reg_9,
	phi_int_arr_reg_8,
	phi_int_arr_reg_7,
	phi_int_arr_reg_6,
	phi_int_arr_reg_5,
	phi_int_arr_reg_4,
	phi_int_arr_reg_3,
	phi_int_arr_reg_2,
	phi_int_arr_reg_1,
	phi_int_arr_reg_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
output 	pipeline_dffe_29;
input 	phi_int_arr_reg_30;
output 	pipeline_dffe_28;
input 	phi_int_arr_reg_31;
input 	phi_int_arr_reg_29;
output 	pipeline_dffe_27;
input 	phi_int_arr_reg_28;
output 	pipeline_dffe_26;
input 	phi_int_arr_reg_27;
output 	pipeline_dffe_25;
input 	phi_int_arr_reg_26;
output 	pipeline_dffe_24;
input 	phi_int_arr_reg_25;
output 	pipeline_dffe_23;
input 	phi_int_arr_reg_24;
output 	pipeline_dffe_22;
input 	phi_int_arr_reg_23;
output 	pipeline_dffe_21;
input 	phi_int_arr_reg_22;
output 	pipeline_dffe_20;
input 	phi_int_arr_reg_21;
output 	pipeline_dffe_19;
input 	phi_int_arr_reg_20;
output 	pipeline_dffe_18;
input 	phi_int_arr_reg_19;
output 	pipeline_dffe_17;
input 	phi_int_arr_reg_18;
output 	pipeline_dffe_16;
input 	phi_int_arr_reg_17;
output 	pipeline_dffe_15;
input 	phi_int_arr_reg_16;
output 	pipeline_dffe_14;
input 	phi_int_arr_reg_15;
output 	pipeline_dffe_13;
input 	phi_int_arr_reg_14;
output 	pipeline_dffe_12;
input 	phi_int_arr_reg_13;
output 	pipeline_dffe_11;
input 	phi_int_arr_reg_12;
input 	phi_int_arr_reg_11;
input 	phi_int_arr_reg_10;
input 	phi_int_arr_reg_9;
input 	phi_int_arr_reg_8;
input 	phi_int_arr_reg_7;
input 	phi_int_arr_reg_6;
input 	phi_int_arr_reg_5;
input 	phi_int_arr_reg_4;
input 	phi_int_arr_reg_3;
input 	phi_int_arr_reg_2;
input 	phi_int_arr_reg_1;
input 	phi_int_arr_reg_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_hth auto_generated(
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_29(pipeline_dffe_29),
	.phi_int_arr_reg_30(phi_int_arr_reg_30),
	.pipeline_dffe_28(pipeline_dffe_28),
	.phi_int_arr_reg_31(phi_int_arr_reg_31),
	.phi_int_arr_reg_29(phi_int_arr_reg_29),
	.pipeline_dffe_27(pipeline_dffe_27),
	.phi_int_arr_reg_28(phi_int_arr_reg_28),
	.pipeline_dffe_26(pipeline_dffe_26),
	.phi_int_arr_reg_27(phi_int_arr_reg_27),
	.pipeline_dffe_25(pipeline_dffe_25),
	.phi_int_arr_reg_26(phi_int_arr_reg_26),
	.pipeline_dffe_24(pipeline_dffe_24),
	.phi_int_arr_reg_25(phi_int_arr_reg_25),
	.pipeline_dffe_23(pipeline_dffe_23),
	.phi_int_arr_reg_24(phi_int_arr_reg_24),
	.pipeline_dffe_22(pipeline_dffe_22),
	.phi_int_arr_reg_23(phi_int_arr_reg_23),
	.pipeline_dffe_21(pipeline_dffe_21),
	.phi_int_arr_reg_22(phi_int_arr_reg_22),
	.pipeline_dffe_20(pipeline_dffe_20),
	.phi_int_arr_reg_21(phi_int_arr_reg_21),
	.pipeline_dffe_19(pipeline_dffe_19),
	.phi_int_arr_reg_20(phi_int_arr_reg_20),
	.pipeline_dffe_18(pipeline_dffe_18),
	.phi_int_arr_reg_19(phi_int_arr_reg_19),
	.pipeline_dffe_17(pipeline_dffe_17),
	.phi_int_arr_reg_18(phi_int_arr_reg_18),
	.pipeline_dffe_16(pipeline_dffe_16),
	.phi_int_arr_reg_17(phi_int_arr_reg_17),
	.pipeline_dffe_15(pipeline_dffe_15),
	.phi_int_arr_reg_16(phi_int_arr_reg_16),
	.pipeline_dffe_14(pipeline_dffe_14),
	.phi_int_arr_reg_15(phi_int_arr_reg_15),
	.pipeline_dffe_13(pipeline_dffe_13),
	.phi_int_arr_reg_14(phi_int_arr_reg_14),
	.pipeline_dffe_12(pipeline_dffe_12),
	.phi_int_arr_reg_13(phi_int_arr_reg_13),
	.pipeline_dffe_11(pipeline_dffe_11),
	.phi_int_arr_reg_12(phi_int_arr_reg_12),
	.phi_int_arr_reg_11(phi_int_arr_reg_11),
	.phi_int_arr_reg_10(phi_int_arr_reg_10),
	.phi_int_arr_reg_9(phi_int_arr_reg_9),
	.phi_int_arr_reg_8(phi_int_arr_reg_8),
	.phi_int_arr_reg_7(phi_int_arr_reg_7),
	.phi_int_arr_reg_6(phi_int_arr_reg_6),
	.phi_int_arr_reg_5(phi_int_arr_reg_5),
	.phi_int_arr_reg_4(phi_int_arr_reg_4),
	.phi_int_arr_reg_3(phi_int_arr_reg_3),
	.phi_int_arr_reg_2(phi_int_arr_reg_2),
	.phi_int_arr_reg_1(phi_int_arr_reg_1),
	.phi_int_arr_reg_0(phi_int_arr_reg_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_hth (
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_29,
	phi_int_arr_reg_30,
	pipeline_dffe_28,
	phi_int_arr_reg_31,
	phi_int_arr_reg_29,
	pipeline_dffe_27,
	phi_int_arr_reg_28,
	pipeline_dffe_26,
	phi_int_arr_reg_27,
	pipeline_dffe_25,
	phi_int_arr_reg_26,
	pipeline_dffe_24,
	phi_int_arr_reg_25,
	pipeline_dffe_23,
	phi_int_arr_reg_24,
	pipeline_dffe_22,
	phi_int_arr_reg_23,
	pipeline_dffe_21,
	phi_int_arr_reg_22,
	pipeline_dffe_20,
	phi_int_arr_reg_21,
	pipeline_dffe_19,
	phi_int_arr_reg_20,
	pipeline_dffe_18,
	phi_int_arr_reg_19,
	pipeline_dffe_17,
	phi_int_arr_reg_18,
	pipeline_dffe_16,
	phi_int_arr_reg_17,
	pipeline_dffe_15,
	phi_int_arr_reg_16,
	pipeline_dffe_14,
	phi_int_arr_reg_15,
	pipeline_dffe_13,
	phi_int_arr_reg_14,
	pipeline_dffe_12,
	phi_int_arr_reg_13,
	pipeline_dffe_11,
	phi_int_arr_reg_12,
	phi_int_arr_reg_11,
	phi_int_arr_reg_10,
	phi_int_arr_reg_9,
	phi_int_arr_reg_8,
	phi_int_arr_reg_7,
	phi_int_arr_reg_6,
	phi_int_arr_reg_5,
	phi_int_arr_reg_4,
	phi_int_arr_reg_3,
	phi_int_arr_reg_2,
	phi_int_arr_reg_1,
	phi_int_arr_reg_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_30;
output 	pipeline_dffe_31;
output 	pipeline_dffe_29;
input 	phi_int_arr_reg_30;
output 	pipeline_dffe_28;
input 	phi_int_arr_reg_31;
input 	phi_int_arr_reg_29;
output 	pipeline_dffe_27;
input 	phi_int_arr_reg_28;
output 	pipeline_dffe_26;
input 	phi_int_arr_reg_27;
output 	pipeline_dffe_25;
input 	phi_int_arr_reg_26;
output 	pipeline_dffe_24;
input 	phi_int_arr_reg_25;
output 	pipeline_dffe_23;
input 	phi_int_arr_reg_24;
output 	pipeline_dffe_22;
input 	phi_int_arr_reg_23;
output 	pipeline_dffe_21;
input 	phi_int_arr_reg_22;
output 	pipeline_dffe_20;
input 	phi_int_arr_reg_21;
output 	pipeline_dffe_19;
input 	phi_int_arr_reg_20;
output 	pipeline_dffe_18;
input 	phi_int_arr_reg_19;
output 	pipeline_dffe_17;
input 	phi_int_arr_reg_18;
output 	pipeline_dffe_16;
input 	phi_int_arr_reg_17;
output 	pipeline_dffe_15;
input 	phi_int_arr_reg_16;
output 	pipeline_dffe_14;
input 	phi_int_arr_reg_15;
output 	pipeline_dffe_13;
input 	phi_int_arr_reg_14;
output 	pipeline_dffe_12;
input 	phi_int_arr_reg_13;
output 	pipeline_dffe_11;
input 	phi_int_arr_reg_12;
input 	phi_int_arr_reg_11;
input 	phi_int_arr_reg_10;
input 	phi_int_arr_reg_9;
input 	phi_int_arr_reg_8;
input 	phi_int_arr_reg_7;
input 	phi_int_arr_reg_6;
input 	phi_int_arr_reg_5;
input 	phi_int_arr_reg_4;
input 	phi_int_arr_reg_3;
input 	phi_int_arr_reg_2;
input 	phi_int_arr_reg_1;
input 	phi_int_arr_reg_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~125_sumout ;
wire \pipeline_dffe[0]~q ;
wire \op_1~126 ;
wire \op_1~121_sumout ;
wire \pipeline_dffe[1]~q ;
wire \op_1~122 ;
wire \op_1~117_sumout ;
wire \pipeline_dffe[2]~q ;
wire \op_1~118 ;
wire \op_1~113_sumout ;
wire \pipeline_dffe[3]~q ;
wire \op_1~114 ;
wire \op_1~109_sumout ;
wire \pipeline_dffe[4]~q ;
wire \op_1~110 ;
wire \op_1~105_sumout ;
wire \pipeline_dffe[5]~q ;
wire \op_1~106 ;
wire \op_1~101_sumout ;
wire \pipeline_dffe[6]~q ;
wire \op_1~102 ;
wire \op_1~97_sumout ;
wire \pipeline_dffe[7]~q ;
wire \op_1~98 ;
wire \op_1~93_sumout ;
wire \pipeline_dffe[8]~q ;
wire \op_1~94 ;
wire \op_1~89_sumout ;
wire \pipeline_dffe[9]~q ;
wire \op_1~90 ;
wire \op_1~85_sumout ;
wire \pipeline_dffe[10]~q ;
wire \op_1~86 ;
wire \op_1~82 ;
wire \op_1~78 ;
wire \op_1~74 ;
wire \op_1~70 ;
wire \op_1~66 ;
wire \op_1~62 ;
wire \op_1~58 ;
wire \op_1~54 ;
wire \op_1~50 ;
wire \op_1~46 ;
wire \op_1~42 ;
wire \op_1~38 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~73_sumout ;
wire \op_1~77_sumout ;
wire \op_1~81_sumout ;


dffeas \pipeline_dffe[30] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_30),
	.prn(vcc));
defparam \pipeline_dffe[30] .is_wysiwyg = "true";
defparam \pipeline_dffe[30] .power_up = "low";

dffeas \pipeline_dffe[31] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_31),
	.prn(vcc));
defparam \pipeline_dffe[31] .is_wysiwyg = "true";
defparam \pipeline_dffe[31] .power_up = "low";

dffeas \pipeline_dffe[29] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_29),
	.prn(vcc));
defparam \pipeline_dffe[29] .is_wysiwyg = "true";
defparam \pipeline_dffe[29] .power_up = "low";

dffeas \pipeline_dffe[28] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_28),
	.prn(vcc));
defparam \pipeline_dffe[28] .is_wysiwyg = "true";
defparam \pipeline_dffe[28] .power_up = "low";

dffeas \pipeline_dffe[27] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_27),
	.prn(vcc));
defparam \pipeline_dffe[27] .is_wysiwyg = "true";
defparam \pipeline_dffe[27] .power_up = "low";

dffeas \pipeline_dffe[26] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_26),
	.prn(vcc));
defparam \pipeline_dffe[26] .is_wysiwyg = "true";
defparam \pipeline_dffe[26] .power_up = "low";

dffeas \pipeline_dffe[25] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_25),
	.prn(vcc));
defparam \pipeline_dffe[25] .is_wysiwyg = "true";
defparam \pipeline_dffe[25] .power_up = "low";

dffeas \pipeline_dffe[24] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_24),
	.prn(vcc));
defparam \pipeline_dffe[24] .is_wysiwyg = "true";
defparam \pipeline_dffe[24] .power_up = "low";

dffeas \pipeline_dffe[23] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_23),
	.prn(vcc));
defparam \pipeline_dffe[23] .is_wysiwyg = "true";
defparam \pipeline_dffe[23] .power_up = "low";

dffeas \pipeline_dffe[22] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_22),
	.prn(vcc));
defparam \pipeline_dffe[22] .is_wysiwyg = "true";
defparam \pipeline_dffe[22] .power_up = "low";

dffeas \pipeline_dffe[21] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_21),
	.prn(vcc));
defparam \pipeline_dffe[21] .is_wysiwyg = "true";
defparam \pipeline_dffe[21] .power_up = "low";

dffeas \pipeline_dffe[20] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \pipeline_dffe[20] .is_wysiwyg = "true";
defparam \pipeline_dffe[20] .power_up = "low";

dffeas \pipeline_dffe[19] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \pipeline_dffe[19] .is_wysiwyg = "true";
defparam \pipeline_dffe[19] .power_up = "low";

dffeas \pipeline_dffe[18] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \pipeline_dffe[18] .is_wysiwyg = "true";
defparam \pipeline_dffe[18] .power_up = "low";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~73_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~77_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~81_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

cyclonev_lcell_comb \op_1~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[0]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~125_sumout ),
	.cout(\op_1~126 ),
	.shareout());
defparam \op_1~125 .extended_lut = "off";
defparam \op_1~125 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~125 .shared_arith = "off";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~125_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[0]~q ),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

cyclonev_lcell_comb \op_1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[1]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_1),
	.datag(gnd),
	.cin(\op_1~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~121_sumout ),
	.cout(\op_1~122 ),
	.shareout());
defparam \op_1~121 .extended_lut = "off";
defparam \op_1~121 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~121 .shared_arith = "off";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~121_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[1]~q ),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

cyclonev_lcell_comb \op_1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[2]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_2),
	.datag(gnd),
	.cin(\op_1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~117_sumout ),
	.cout(\op_1~118 ),
	.shareout());
defparam \op_1~117 .extended_lut = "off";
defparam \op_1~117 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~117 .shared_arith = "off";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~117_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[2]~q ),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

cyclonev_lcell_comb \op_1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[3]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_3),
	.datag(gnd),
	.cin(\op_1~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~113_sumout ),
	.cout(\op_1~114 ),
	.shareout());
defparam \op_1~113 .extended_lut = "off";
defparam \op_1~113 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~113 .shared_arith = "off";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~113_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[3]~q ),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

cyclonev_lcell_comb \op_1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[4]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_4),
	.datag(gnd),
	.cin(\op_1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~109_sumout ),
	.cout(\op_1~110 ),
	.shareout());
defparam \op_1~109 .extended_lut = "off";
defparam \op_1~109 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~109 .shared_arith = "off";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~109_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[4]~q ),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

cyclonev_lcell_comb \op_1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[5]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_5),
	.datag(gnd),
	.cin(\op_1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~105_sumout ),
	.cout(\op_1~106 ),
	.shareout());
defparam \op_1~105 .extended_lut = "off";
defparam \op_1~105 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~105 .shared_arith = "off";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~105_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[5]~q ),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

cyclonev_lcell_comb \op_1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[6]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_6),
	.datag(gnd),
	.cin(\op_1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~101_sumout ),
	.cout(\op_1~102 ),
	.shareout());
defparam \op_1~101 .extended_lut = "off";
defparam \op_1~101 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~101 .shared_arith = "off";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~101_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[6]~q ),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

cyclonev_lcell_comb \op_1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[7]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_7),
	.datag(gnd),
	.cin(\op_1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~97_sumout ),
	.cout(\op_1~98 ),
	.shareout());
defparam \op_1~97 .extended_lut = "off";
defparam \op_1~97 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~97 .shared_arith = "off";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~97_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[7]~q ),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

cyclonev_lcell_comb \op_1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[8]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_8),
	.datag(gnd),
	.cin(\op_1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~93_sumout ),
	.cout(\op_1~94 ),
	.shareout());
defparam \op_1~93 .extended_lut = "off";
defparam \op_1~93 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~93 .shared_arith = "off";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~93_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[8]~q ),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

cyclonev_lcell_comb \op_1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[9]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_9),
	.datag(gnd),
	.cin(\op_1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~89_sumout ),
	.cout(\op_1~90 ),
	.shareout());
defparam \op_1~89 .extended_lut = "off";
defparam \op_1~89 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~89 .shared_arith = "off";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~89_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[9]~q ),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \op_1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\pipeline_dffe[10]~q ),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_10),
	.datag(gnd),
	.cin(\op_1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~85_sumout ),
	.cout(\op_1~86 ),
	.shareout());
defparam \op_1~85 .extended_lut = "off";
defparam \op_1~85 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~85 .shared_arith = "off";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~85_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[10]~q ),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

cyclonev_lcell_comb \op_1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_11),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_11),
	.datag(gnd),
	.cin(\op_1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~81_sumout ),
	.cout(\op_1~82 ),
	.shareout());
defparam \op_1~81 .extended_lut = "off";
defparam \op_1~81 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~81 .shared_arith = "off";

cyclonev_lcell_comb \op_1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_12),
	.datag(gnd),
	.cin(\op_1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~77_sumout ),
	.cout(\op_1~78 ),
	.shareout());
defparam \op_1~77 .extended_lut = "off";
defparam \op_1~77 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~77 .shared_arith = "off";

cyclonev_lcell_comb \op_1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_13),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_13),
	.datag(gnd),
	.cin(\op_1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~73_sumout ),
	.cout(\op_1~74 ),
	.shareout());
defparam \op_1~73 .extended_lut = "off";
defparam \op_1~73 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~73 .shared_arith = "off";

cyclonev_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_14),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_14),
	.datag(gnd),
	.cin(\op_1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

cyclonev_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_15),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_15),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

cyclonev_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_16),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_16),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

cyclonev_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_17),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_17),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

cyclonev_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_18),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

cyclonev_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_19),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_19),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_20),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_20),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_21),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_22),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_22),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_23),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_23),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_24),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_24),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_25),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_25),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_26),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_26),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_27),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_27),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_28),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_28),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_29),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_29),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_30),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_30),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(!phi_int_arr_reg_31),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

endmodule

module NCO_Lab3_asj_crs_par (
	ram_block8a1,
	ram_block8a0,
	sin_o_0,
	sin_o_1,
	sin_o_2,
	sin_o_3,
	sin_o_4,
	sin_o_5,
	sin_o_6,
	sin_o_7,
	sin_o_8,
	sin_o_9,
	sin_o_10,
	sin_o_11,
	cordic_x_res_2c_0,
	cordic_y_res_2c_0,
	cordic_y_res_d_1,
	cordic_x_res_d_1,
	cordic_y_res_2c_1,
	cordic_x_res_2c_1,
	cordic_y_res_d_2,
	cordic_x_res_d_2,
	cordic_y_res_2c_2,
	cordic_x_res_2c_2,
	cordic_y_res_d_3,
	cordic_x_res_d_3,
	cordic_y_res_2c_3,
	cordic_x_res_2c_3,
	cordic_y_res_d_4,
	cordic_x_res_d_4,
	cordic_y_res_2c_4,
	cordic_x_res_2c_4,
	cordic_y_res_d_5,
	cordic_x_res_d_5,
	cordic_y_res_2c_5,
	cordic_x_res_2c_5,
	cordic_y_res_d_6,
	cordic_x_res_d_6,
	cordic_y_res_2c_6,
	cordic_x_res_2c_6,
	cordic_y_res_d_7,
	cordic_x_res_d_7,
	cordic_y_res_2c_7,
	cordic_x_res_2c_7,
	cordic_y_res_d_8,
	cordic_x_res_d_8,
	cordic_y_res_2c_8,
	cordic_x_res_2c_8,
	cordic_y_res_d_9,
	cordic_x_res_d_9,
	cordic_y_res_2c_9,
	cordic_x_res_2c_9,
	cordic_y_res_d_10,
	cordic_x_res_d_10,
	cordic_y_res_2c_10,
	cordic_x_res_2c_10,
	cordic_y_res_d_11,
	cordic_x_res_d_11,
	cordic_y_res_2c_11,
	cordic_x_res_2c_11,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	ram_block8a1;
input 	ram_block8a0;
output 	sin_o_0;
output 	sin_o_1;
output 	sin_o_2;
output 	sin_o_3;
output 	sin_o_4;
output 	sin_o_5;
output 	sin_o_6;
output 	sin_o_7;
output 	sin_o_8;
output 	sin_o_9;
output 	sin_o_10;
output 	sin_o_11;
input 	cordic_x_res_2c_0;
input 	cordic_y_res_2c_0;
input 	cordic_y_res_d_1;
input 	cordic_x_res_d_1;
input 	cordic_y_res_2c_1;
input 	cordic_x_res_2c_1;
input 	cordic_y_res_d_2;
input 	cordic_x_res_d_2;
input 	cordic_y_res_2c_2;
input 	cordic_x_res_2c_2;
input 	cordic_y_res_d_3;
input 	cordic_x_res_d_3;
input 	cordic_y_res_2c_3;
input 	cordic_x_res_2c_3;
input 	cordic_y_res_d_4;
input 	cordic_x_res_d_4;
input 	cordic_y_res_2c_4;
input 	cordic_x_res_2c_4;
input 	cordic_y_res_d_5;
input 	cordic_x_res_d_5;
input 	cordic_y_res_2c_5;
input 	cordic_x_res_2c_5;
input 	cordic_y_res_d_6;
input 	cordic_x_res_d_6;
input 	cordic_y_res_2c_6;
input 	cordic_x_res_2c_6;
input 	cordic_y_res_d_7;
input 	cordic_x_res_d_7;
input 	cordic_y_res_2c_7;
input 	cordic_x_res_2c_7;
input 	cordic_y_res_d_8;
input 	cordic_x_res_d_8;
input 	cordic_y_res_2c_8;
input 	cordic_x_res_2c_8;
input 	cordic_y_res_d_9;
input 	cordic_x_res_d_9;
input 	cordic_y_res_2c_9;
input 	cordic_x_res_2c_9;
input 	cordic_y_res_d_10;
input 	cordic_x_res_d_10;
input 	cordic_y_res_2c_10;
input 	cordic_x_res_2c_10;
input 	cordic_y_res_d_11;
input 	cordic_x_res_d_11;
input 	cordic_y_res_2c_11;
input 	cordic_x_res_2c_11;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Mux11~0_combout ;
wire \Mux10~0_combout ;
wire \Mux9~0_combout ;
wire \Mux8~0_combout ;
wire \Mux7~0_combout ;
wire \Mux6~0_combout ;
wire \Mux5~0_combout ;
wire \Mux4~0_combout ;
wire \Mux3~0_combout ;
wire \Mux2~0_combout ;
wire \Mux1~0_combout ;
wire \Mux0~0_combout ;


dffeas \sin_o[0] (
	.clk(clk),
	.d(\Mux11~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_0),
	.prn(vcc));
defparam \sin_o[0] .is_wysiwyg = "true";
defparam \sin_o[0] .power_up = "low";

dffeas \sin_o[1] (
	.clk(clk),
	.d(\Mux10~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_1),
	.prn(vcc));
defparam \sin_o[1] .is_wysiwyg = "true";
defparam \sin_o[1] .power_up = "low";

dffeas \sin_o[2] (
	.clk(clk),
	.d(\Mux9~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_2),
	.prn(vcc));
defparam \sin_o[2] .is_wysiwyg = "true";
defparam \sin_o[2] .power_up = "low";

dffeas \sin_o[3] (
	.clk(clk),
	.d(\Mux8~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_3),
	.prn(vcc));
defparam \sin_o[3] .is_wysiwyg = "true";
defparam \sin_o[3] .power_up = "low";

dffeas \sin_o[4] (
	.clk(clk),
	.d(\Mux7~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_4),
	.prn(vcc));
defparam \sin_o[4] .is_wysiwyg = "true";
defparam \sin_o[4] .power_up = "low";

dffeas \sin_o[5] (
	.clk(clk),
	.d(\Mux6~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_5),
	.prn(vcc));
defparam \sin_o[5] .is_wysiwyg = "true";
defparam \sin_o[5] .power_up = "low";

dffeas \sin_o[6] (
	.clk(clk),
	.d(\Mux5~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_6),
	.prn(vcc));
defparam \sin_o[6] .is_wysiwyg = "true";
defparam \sin_o[6] .power_up = "low";

dffeas \sin_o[7] (
	.clk(clk),
	.d(\Mux4~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_7),
	.prn(vcc));
defparam \sin_o[7] .is_wysiwyg = "true";
defparam \sin_o[7] .power_up = "low";

dffeas \sin_o[8] (
	.clk(clk),
	.d(\Mux3~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_8),
	.prn(vcc));
defparam \sin_o[8] .is_wysiwyg = "true";
defparam \sin_o[8] .power_up = "low";

dffeas \sin_o[9] (
	.clk(clk),
	.d(\Mux2~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_9),
	.prn(vcc));
defparam \sin_o[9] .is_wysiwyg = "true";
defparam \sin_o[9] .power_up = "low";

dffeas \sin_o[10] (
	.clk(clk),
	.d(\Mux1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_10),
	.prn(vcc));
defparam \sin_o[10] .is_wysiwyg = "true";
defparam \sin_o[10] .power_up = "low";

dffeas \sin_o[11] (
	.clk(clk),
	.d(\Mux0~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_11),
	.prn(vcc));
defparam \sin_o[11] .is_wysiwyg = "true";
defparam \sin_o[11] .power_up = "low";

cyclonev_lcell_comb \Mux11~0 (
	.dataa(!cordic_x_res_2c_0),
	.datab(!ram_block8a1),
	.datac(!cordic_y_res_2c_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux11~0 .extended_lut = "off";
defparam \Mux11~0 .lut_mask = 64'h4747474747474747;
defparam \Mux11~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux10~0 (
	.dataa(!cordic_y_res_d_1),
	.datab(!cordic_x_res_d_1),
	.datac(!cordic_y_res_2c_1),
	.datad(!cordic_x_res_2c_1),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux10~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux10~0 .extended_lut = "off";
defparam \Mux10~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux10~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux9~0 (
	.dataa(!cordic_y_res_d_2),
	.datab(!cordic_x_res_d_2),
	.datac(!cordic_y_res_2c_2),
	.datad(!cordic_x_res_2c_2),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux9~0 .extended_lut = "off";
defparam \Mux9~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux9~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux8~0 (
	.dataa(!cordic_y_res_d_3),
	.datab(!cordic_x_res_d_3),
	.datac(!cordic_y_res_2c_3),
	.datad(!cordic_x_res_2c_3),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux8~0 .extended_lut = "off";
defparam \Mux8~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux8~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux7~0 (
	.dataa(!cordic_y_res_d_4),
	.datab(!cordic_x_res_d_4),
	.datac(!cordic_y_res_2c_4),
	.datad(!cordic_x_res_2c_4),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux7~0 .extended_lut = "off";
defparam \Mux7~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux7~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux6~0 (
	.dataa(!cordic_y_res_d_5),
	.datab(!cordic_x_res_d_5),
	.datac(!cordic_y_res_2c_5),
	.datad(!cordic_x_res_2c_5),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux6~0 .extended_lut = "off";
defparam \Mux6~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux6~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux5~0 (
	.dataa(!cordic_y_res_d_6),
	.datab(!cordic_x_res_d_6),
	.datac(!cordic_y_res_2c_6),
	.datad(!cordic_x_res_2c_6),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux5~0 .extended_lut = "off";
defparam \Mux5~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux5~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux4~0 (
	.dataa(!cordic_y_res_d_7),
	.datab(!cordic_x_res_d_7),
	.datac(!cordic_y_res_2c_7),
	.datad(!cordic_x_res_2c_7),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux4~0 .extended_lut = "off";
defparam \Mux4~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux4~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux3~0 (
	.dataa(!cordic_y_res_d_8),
	.datab(!cordic_x_res_d_8),
	.datac(!cordic_y_res_2c_8),
	.datad(!cordic_x_res_2c_8),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux3~0 .extended_lut = "off";
defparam \Mux3~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux3~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!cordic_y_res_d_9),
	.datab(!cordic_x_res_d_9),
	.datac(!cordic_y_res_2c_9),
	.datad(!cordic_x_res_2c_9),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux1~0 (
	.dataa(!cordic_y_res_d_10),
	.datab(!cordic_x_res_d_10),
	.datac(!cordic_y_res_2c_10),
	.datad(!cordic_x_res_2c_10),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux1~0 .extended_lut = "off";
defparam \Mux1~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux1~0 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!cordic_y_res_d_11),
	.datab(!cordic_x_res_d_11),
	.datac(!cordic_y_res_2c_11),
	.datad(!cordic_x_res_2c_11),
	.datae(!ram_block8a1),
	.dataf(!ram_block8a0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "off";
defparam \Mux0~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux0~0 .shared_arith = "off";

endmodule

module NCO_Lab3_asj_dxx (
	ram_block8a1,
	ram_block8a0,
	dxxrv_3,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_20,
	pipeline_dffe_19,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	dxxrv_2,
	pipeline_dffe_13,
	dxxrv_1,
	pipeline_dffe_12,
	dxxrv_0,
	pipeline_dffe_11,
	dxxpdo_18,
	dxxpdo_17,
	dxxpdo_16,
	dxxpdo_15,
	dxxpdo_14,
	dxxpdo_13,
	dxxpdo_12,
	dxxpdo_11,
	dxxpdo_10,
	dxxpdo_9,
	dxxpdo_8,
	dxxpdo_7,
	dxxpdo_6,
	dxxpdo_5,
	dxxpdo_4,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	ram_block8a1;
output 	ram_block8a0;
input 	dxxrv_3;
input 	pipeline_dffe_30;
input 	pipeline_dffe_31;
input 	pipeline_dffe_29;
input 	pipeline_dffe_28;
input 	pipeline_dffe_27;
input 	pipeline_dffe_26;
input 	pipeline_dffe_25;
input 	pipeline_dffe_24;
input 	pipeline_dffe_23;
input 	pipeline_dffe_22;
input 	pipeline_dffe_21;
input 	pipeline_dffe_20;
input 	pipeline_dffe_19;
input 	pipeline_dffe_18;
input 	pipeline_dffe_17;
input 	pipeline_dffe_16;
input 	pipeline_dffe_15;
input 	pipeline_dffe_14;
input 	dxxrv_2;
input 	pipeline_dffe_13;
input 	dxxrv_1;
input 	pipeline_dffe_12;
input 	dxxrv_0;
input 	pipeline_dffe_11;
output 	dxxpdo_18;
output 	dxxpdo_17;
output 	dxxpdo_16;
output 	dxxpdo_15;
output 	dxxpdo_14;
output 	dxxpdo_13;
output 	dxxpdo_12;
output 	dxxpdo_11;
output 	dxxpdo_10;
output 	dxxpdo_9;
output 	dxxpdo_8;
output 	dxxpdo_7;
output 	dxxpdo_6;
output 	dxxpdo_5;
output 	dxxpdo_4;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ux014|auto_generated|pipeline_dffe[19]~q ;
wire \ux014|auto_generated|pipeline_dffe[20]~q ;
wire \ux014|auto_generated|pipeline_dffe[18]~q ;
wire \ux014|auto_generated|pipeline_dffe[17]~q ;
wire \ux014|auto_generated|pipeline_dffe[16]~q ;
wire \ux014|auto_generated|pipeline_dffe[15]~q ;
wire \ux014|auto_generated|pipeline_dffe[14]~q ;
wire \ux014|auto_generated|pipeline_dffe[13]~q ;
wire \ux014|auto_generated|pipeline_dffe[12]~q ;
wire \ux014|auto_generated|pipeline_dffe[11]~q ;
wire \ux014|auto_generated|pipeline_dffe[10]~q ;
wire \ux014|auto_generated|pipeline_dffe[9]~q ;
wire \ux014|auto_generated|pipeline_dffe[8]~q ;
wire \ux014|auto_generated|pipeline_dffe[7]~q ;
wire \ux014|auto_generated|pipeline_dffe[6]~q ;
wire \ux014|auto_generated|pipeline_dffe[5]~q ;
wire \ux014|auto_generated|pipeline_dffe[4]~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~1_combout ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ;
wire \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~1_sumout ;
wire \dxxpdo_rtl_0|auto_generated|dffe7~0_combout ;
wire \dxxpdo_rtl_0|auto_generated|dffe7~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~1_sumout ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|cout_actual~combout ;
wire \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ;
wire \dxxpdo_rtl_0|auto_generated|op_2~0_combout ;
wire \dxxpdo_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ;
wire \dxxpdo_rtl_0|auto_generated|op_1~1_sumout ;
wire \dxxpdo_rtl_0|auto_generated|dffe3a[0]~q ;
wire \dxxpdo_rtl_0|auto_generated|op_1~2 ;
wire \dxxpdo_rtl_0|auto_generated|op_1~5_sumout ;
wire \dxxpdo_rtl_0|auto_generated|dffe3a[1]~0_combout ;
wire \dxxpdo_rtl_0|auto_generated|dffe3a[1]~q ;
wire \dxxpdo_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ;
wire \dxxpdo_rtl_0|auto_generated|op_1~6 ;
wire \dxxpdo_rtl_0|auto_generated|op_1~9_sumout ;
wire \dxxpdo_rtl_0|auto_generated|dffe3a[2]~q ;
wire \dxxpdo_rtl_0|auto_generated|op_1~10 ;
wire \dxxpdo_rtl_0|auto_generated|op_1~13_sumout ;
wire \dxxpdo_rtl_0|auto_generated|dffe3a[3]~q ;
wire \dxxpdo_rtl_0|auto_generated|op_1~14 ;
wire \dxxpdo_rtl_0|auto_generated|op_1~17_sumout ;
wire \dxxpdo_rtl_0|auto_generated|dffe3a[4]~q ;

wire [143:0] \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1_PORTBDATAOUT_bus ;
wire [143:0] \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus ;

assign ram_block8a1 = \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1_PORTBDATAOUT_bus [0];

assign ram_block8a0 = \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus [0];

NCO_Lab3_lpm_add_sub_2 ux014(
	.pipeline_dffe_19(\ux014|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_20(\ux014|auto_generated|pipeline_dffe[20]~q ),
	.dxxrv_3(dxxrv_3),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_201(pipeline_dffe_20),
	.pipeline_dffe_191(pipeline_dffe_19),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.dxxrv_2(dxxrv_2),
	.pipeline_dffe_13(pipeline_dffe_13),
	.dxxrv_1(dxxrv_1),
	.pipeline_dffe_12(pipeline_dffe_12),
	.dxxrv_0(dxxrv_0),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_181(\ux014|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_171(\ux014|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_161(\ux014|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_151(\ux014|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_141(\ux014|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_131(\ux014|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_121(\ux014|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_111(\ux014|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\ux014|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\ux014|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\ux014|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\ux014|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\ux014|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\ux014|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\ux014|auto_generated|pipeline_dffe[4]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_ram_block \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(clken),
	.ena1(clken),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\dxxpdo_rtl_0|auto_generated|dffe7~q ),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\ux014|auto_generated|pipeline_dffe[19]~q }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,
\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\dxxpdo_rtl_0|auto_generated|dffe3a[4]~q ,\dxxpdo_rtl_0|auto_generated|dffe3a[3]~q ,\dxxpdo_rtl_0|auto_generated|dffe3a[2]~q ,\dxxpdo_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\dxxpdo_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .clk0_core_clock_enable = "ena0";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .clk0_input_clock_enable = "ena0";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .clk1_output_clock_enable = "ena1";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .data_interleave_offset_in_bits = 1;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .data_interleave_width_in_bits = 1;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .logical_ram_name = "NCO_Lab3_nco_ii_0:nco_ii_0|asj_dxx:ux002|altshift_taps:dxxpdo_rtl_0|shift_taps_duv:auto_generated|altsyncram_pfc1:altsyncram5|ALTSYNCRAM";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .mixed_port_feed_through_mode = "dont_care";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .operation_mode = "dual_port";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_address_clear = "none";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_address_width = 5;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_data_out_clear = "none";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_data_out_clock = "none";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_data_width = 1;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_first_address = 0;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_first_bit_number = 1;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_last_address = 26;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_logical_ram_depth = 27;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_logical_ram_width = 2;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_address_clear = "none";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_address_clock = "clock0";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_address_width = 5;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_data_out_clear = "clear0";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_data_out_clock = "clock1";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_data_width = 1;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_first_address = 0;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_first_bit_number = 1;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_last_address = 26;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_logical_ram_depth = 27;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_logical_ram_width = 2;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .port_b_read_enable_clock = "clock0";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a1 .ram_block_type = "auto";

cyclonev_ram_block \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 (
	.portawe(vcc),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(clk),
	.ena0(clken),
	.ena1(clken),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!\dxxpdo_rtl_0|auto_generated|dffe7~q ),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\ux014|auto_generated|pipeline_dffe[20]~q }),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ,\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ,\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ,
\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ,\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\dxxpdo_rtl_0|auto_generated|dffe3a[4]~q ,\dxxpdo_rtl_0|auto_generated|dffe3a[3]~q ,\dxxpdo_rtl_0|auto_generated|dffe3a[2]~q ,\dxxpdo_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ,\dxxpdo_rtl_0|auto_generated|dffe3a[0]~q }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0_PORTBDATAOUT_bus ),
	.eccstatus(),
	.dftout());
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk0_core_clock_enable = "ena0";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk0_input_clock_enable = "ena0";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .clk1_output_clock_enable = "ena1";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .data_interleave_offset_in_bits = 1;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .data_interleave_width_in_bits = 1;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .logical_ram_name = "NCO_Lab3_nco_ii_0:nco_ii_0|asj_dxx:ux002|altshift_taps:dxxpdo_rtl_0|shift_taps_duv:auto_generated|altsyncram_pfc1:altsyncram5|ALTSYNCRAM";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .mixed_port_feed_through_mode = "dont_care";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .operation_mode = "dual_port";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_address_clear = "none";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_address_width = 5;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_out_clear = "none";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_out_clock = "none";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_data_width = 1;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_first_address = 0;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_first_bit_number = 0;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_last_address = 26;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_logical_ram_depth = 27;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_logical_ram_width = 2;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_clear = "none";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_clock = "clock0";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_address_width = 5;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_out_clear = "clear0";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_out_clock = "clock1";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_data_width = 1;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_first_address = 0;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_first_bit_number = 0;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_last_address = 26;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_logical_ram_depth = 27;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_logical_ram_width = 2;
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .port_b_read_enable_clock = "clock0";
defparam \dxxpdo_rtl_0|auto_generated|altsyncram5|ram_block8a0 .ram_block_type = "auto";

dffeas \dxxpdo[18] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[18]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_18),
	.prn(vcc));
defparam \dxxpdo[18] .is_wysiwyg = "true";
defparam \dxxpdo[18] .power_up = "low";

dffeas \dxxpdo[17] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[17]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_17),
	.prn(vcc));
defparam \dxxpdo[17] .is_wysiwyg = "true";
defparam \dxxpdo[17] .power_up = "low";

dffeas \dxxpdo[16] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[16]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_16),
	.prn(vcc));
defparam \dxxpdo[16] .is_wysiwyg = "true";
defparam \dxxpdo[16] .power_up = "low";

dffeas \dxxpdo[15] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[15]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_15),
	.prn(vcc));
defparam \dxxpdo[15] .is_wysiwyg = "true";
defparam \dxxpdo[15] .power_up = "low";

dffeas \dxxpdo[14] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[14]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_14),
	.prn(vcc));
defparam \dxxpdo[14] .is_wysiwyg = "true";
defparam \dxxpdo[14] .power_up = "low";

dffeas \dxxpdo[13] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[13]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_13),
	.prn(vcc));
defparam \dxxpdo[13] .is_wysiwyg = "true";
defparam \dxxpdo[13] .power_up = "low";

dffeas \dxxpdo[12] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[12]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_12),
	.prn(vcc));
defparam \dxxpdo[12] .is_wysiwyg = "true";
defparam \dxxpdo[12] .power_up = "low";

dffeas \dxxpdo[11] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[11]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_11),
	.prn(vcc));
defparam \dxxpdo[11] .is_wysiwyg = "true";
defparam \dxxpdo[11] .power_up = "low";

dffeas \dxxpdo[10] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[10]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_10),
	.prn(vcc));
defparam \dxxpdo[10] .is_wysiwyg = "true";
defparam \dxxpdo[10] .power_up = "low";

dffeas \dxxpdo[9] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_9),
	.prn(vcc));
defparam \dxxpdo[9] .is_wysiwyg = "true";
defparam \dxxpdo[9] .power_up = "low";

dffeas \dxxpdo[8] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_8),
	.prn(vcc));
defparam \dxxpdo[8] .is_wysiwyg = "true";
defparam \dxxpdo[8] .power_up = "low";

dffeas \dxxpdo[7] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[7]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_7),
	.prn(vcc));
defparam \dxxpdo[7] .is_wysiwyg = "true";
defparam \dxxpdo[7] .power_up = "low";

dffeas \dxxpdo[6] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[6]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_6),
	.prn(vcc));
defparam \dxxpdo[6] .is_wysiwyg = "true";
defparam \dxxpdo[6] .power_up = "low";

dffeas \dxxpdo[5] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[5]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_5),
	.prn(vcc));
defparam \dxxpdo[5] .is_wysiwyg = "true";
defparam \dxxpdo[5] .power_up = "low";

dffeas \dxxpdo[4] (
	.clk(clk),
	.d(\ux014|auto_generated|pipeline_dffe[4]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxpdo_4),
	.prn(vcc));
defparam \dxxpdo[4] .is_wysiwyg = "true";
defparam \dxxpdo[4] .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita0 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita0 .lut_mask = 64'h000000000000FF00;
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita0 .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 (
	.dataa(!\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita0~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~1 .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 (
	.dataa(!clken),
	.datab(!\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~1_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .lut_mask = 64'h7777777777777777;
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0 (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0 .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0 .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita1 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita1 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit1 (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit1~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit1 .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit1 .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita2 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita2 .lut_mask = 64'h00000000000000FF;
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita2 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit2 (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit2~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit2 .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit2 .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita3 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita3 .lut_mask = 64'h000000000000FF00;
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita3 .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 (
	.dataa(!\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita3~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3~0 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3 (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3 .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit3 .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4 .lut_mask = 64'h000000000000FF00;
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4 .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 (
	.dataa(!\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4~0 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4 (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit0~0_combout ),
	.q(\dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4 .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_reg_bit4 .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~1_sumout ),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~1 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~1 .lut_mask = 64'h0000000000000000;
defparam \dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~1 .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|dffe7~0 (
	.dataa(!\dxxpdo_rtl_0|auto_generated|cntr6|counter_comb_bita4~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dxxpdo_rtl_0|auto_generated|dffe7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|dffe7~0 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|dffe7~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dxxpdo_rtl_0|auto_generated|dffe7~0 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|dffe7 (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|dffe7~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|dffe7~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|dffe7 .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|dffe7 .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita0 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita0 .lut_mask = 64'h00000000000000FF;
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita0 .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita1 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita1 .lut_mask = 64'h00000000000000FF;
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita1 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1] (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dxxpdo_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1] .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita2 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita2 .lut_mask = 64'h00000000000000FF;
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita2 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2] (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dxxpdo_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita3 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita3 .lut_mask = 64'h00000000000000FF;
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita3 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3] (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dxxpdo_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3] .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4 .lut_mask = 64'h00000000000000FF;
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4] (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dxxpdo_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4] .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~1_sumout ),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 .lut_mask = 64'h0000000000000000;
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~1 .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cntr1|cout_actual (
	.dataa(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.dataf(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita4~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dxxpdo_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cntr1|cout_actual .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|cout_actual .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \dxxpdo_rtl_0|auto_generated|cntr1|cout_actual .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0] (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|cntr1|counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\dxxpdo_rtl_0|auto_generated|cntr1|cout_actual~combout ),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0] .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|op_2~0 (
	.dataa(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dxxpdo_rtl_0|auto_generated|op_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|op_2~0 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|op_2~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \dxxpdo_rtl_0|auto_generated|op_2~0 .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|cmpr4_aeb_int~0 (
	.dataa(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datab(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datac(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dxxpdo_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|cmpr4_aeb_int~0 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|cmpr4_aeb_int~0 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \dxxpdo_rtl_0|auto_generated|cmpr4_aeb_int~0 .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|op_1~1 (
	.dataa(!\dxxpdo_rtl_0|auto_generated|op_2~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[0]~q ),
	.datae(gnd),
	.dataf(!\dxxpdo_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|op_1~1_sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|op_1~2 ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|op_1~1 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|op_1~1 .lut_mask = 64'h000055FF000000FF;
defparam \dxxpdo_rtl_0|auto_generated|op_1~1 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|dffe3a[0] (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|op_1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|dffe3a[0]~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[0] .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[0] .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|op_1~5 (
	.dataa(!\dxxpdo_rtl_0|auto_generated|op_2~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[1]~q ),
	.datae(gnd),
	.dataf(!\dxxpdo_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|op_1~5_sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|op_1~6 ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|op_1~5 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|op_1~5 .lut_mask = 64'h000055FF000000FF;
defparam \dxxpdo_rtl_0|auto_generated|op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|dffe3a[1]~0 (
	.dataa(!\dxxpdo_rtl_0|auto_generated|op_1~5_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dxxpdo_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[1]~0 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[1]~0 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|dffe3a[1] (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|dffe3a[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|dffe3a[1]~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[1] .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[1] .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|dffe3a[1]~_wirecell (
	.dataa(!\dxxpdo_rtl_0|auto_generated|dffe3a[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dxxpdo_rtl_0|auto_generated|dffe3a[1]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[1]~_wirecell .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[1]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[1]~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|op_1~9_sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|op_1~10 ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|op_1~9 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|op_1~9 .lut_mask = 64'h00000000000000FF;
defparam \dxxpdo_rtl_0|auto_generated|op_1~9 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|dffe3a[2] (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|op_1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|dffe3a[2]~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[2] .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[2] .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|op_1~13 (
	.dataa(!\dxxpdo_rtl_0|auto_generated|op_2~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(!\dxxpdo_rtl_0|auto_generated|cmpr4_aeb_int~0_combout ),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|op_1~13_sumout ),
	.cout(\dxxpdo_rtl_0|auto_generated|op_1~14 ),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|op_1~13 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|op_1~13 .lut_mask = 64'h0000FFAA000000FF;
defparam \dxxpdo_rtl_0|auto_generated|op_1~13 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|dffe3a[3] (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|op_1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|dffe3a[3]~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[3] .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[3] .power_up = "low";

cyclonev_lcell_comb \dxxpdo_rtl_0|auto_generated|op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\dxxpdo_rtl_0|auto_generated|cntr1|counter_reg_bit[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\dxxpdo_rtl_0|auto_generated|op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\dxxpdo_rtl_0|auto_generated|op_1~17_sumout ),
	.cout(),
	.shareout());
defparam \dxxpdo_rtl_0|auto_generated|op_1~17 .extended_lut = "off";
defparam \dxxpdo_rtl_0|auto_generated|op_1~17 .lut_mask = 64'h00000000000000FF;
defparam \dxxpdo_rtl_0|auto_generated|op_1~17 .shared_arith = "off";

dffeas \dxxpdo_rtl_0|auto_generated|dffe3a[4] (
	.clk(clk),
	.d(\dxxpdo_rtl_0|auto_generated|op_1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\dxxpdo_rtl_0|auto_generated|dffe3a[4]~q ),
	.prn(vcc));
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[4] .is_wysiwyg = "true";
defparam \dxxpdo_rtl_0|auto_generated|dffe3a[4] .power_up = "low";

endmodule

module NCO_Lab3_lpm_add_sub_2 (
	pipeline_dffe_19,
	pipeline_dffe_20,
	dxxrv_3,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_201,
	pipeline_dffe_191,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	dxxrv_2,
	pipeline_dffe_13,
	dxxrv_1,
	pipeline_dffe_12,
	dxxrv_0,
	pipeline_dffe_11,
	pipeline_dffe_181,
	pipeline_dffe_171,
	pipeline_dffe_161,
	pipeline_dffe_151,
	pipeline_dffe_141,
	pipeline_dffe_131,
	pipeline_dffe_121,
	pipeline_dffe_111,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
input 	dxxrv_3;
input 	pipeline_dffe_30;
input 	pipeline_dffe_31;
input 	pipeline_dffe_29;
input 	pipeline_dffe_28;
input 	pipeline_dffe_27;
input 	pipeline_dffe_26;
input 	pipeline_dffe_25;
input 	pipeline_dffe_24;
input 	pipeline_dffe_23;
input 	pipeline_dffe_22;
input 	pipeline_dffe_21;
input 	pipeline_dffe_201;
input 	pipeline_dffe_191;
input 	pipeline_dffe_18;
input 	pipeline_dffe_17;
input 	pipeline_dffe_16;
input 	pipeline_dffe_15;
input 	pipeline_dffe_14;
input 	dxxrv_2;
input 	pipeline_dffe_13;
input 	dxxrv_1;
input 	pipeline_dffe_12;
input 	dxxrv_0;
input 	pipeline_dffe_11;
output 	pipeline_dffe_181;
output 	pipeline_dffe_171;
output 	pipeline_dffe_161;
output 	pipeline_dffe_151;
output 	pipeline_dffe_141;
output 	pipeline_dffe_131;
output 	pipeline_dffe_121;
output 	pipeline_dffe_111;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_cmh auto_generated(
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_20(pipeline_dffe_20),
	.dxxrv_3(dxxrv_3),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_201(pipeline_dffe_201),
	.pipeline_dffe_191(pipeline_dffe_191),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.dxxrv_2(dxxrv_2),
	.pipeline_dffe_13(pipeline_dffe_13),
	.dxxrv_1(dxxrv_1),
	.pipeline_dffe_12(pipeline_dffe_12),
	.dxxrv_0(dxxrv_0),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_181(pipeline_dffe_181),
	.pipeline_dffe_171(pipeline_dffe_171),
	.pipeline_dffe_161(pipeline_dffe_161),
	.pipeline_dffe_151(pipeline_dffe_151),
	.pipeline_dffe_141(pipeline_dffe_141),
	.pipeline_dffe_131(pipeline_dffe_131),
	.pipeline_dffe_121(pipeline_dffe_121),
	.pipeline_dffe_111(pipeline_dffe_111),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_cmh (
	pipeline_dffe_19,
	pipeline_dffe_20,
	dxxrv_3,
	pipeline_dffe_30,
	pipeline_dffe_31,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_201,
	pipeline_dffe_191,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	dxxrv_2,
	pipeline_dffe_13,
	dxxrv_1,
	pipeline_dffe_12,
	dxxrv_0,
	pipeline_dffe_11,
	pipeline_dffe_181,
	pipeline_dffe_171,
	pipeline_dffe_161,
	pipeline_dffe_151,
	pipeline_dffe_141,
	pipeline_dffe_131,
	pipeline_dffe_121,
	pipeline_dffe_111,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_19;
output 	pipeline_dffe_20;
input 	dxxrv_3;
input 	pipeline_dffe_30;
input 	pipeline_dffe_31;
input 	pipeline_dffe_29;
input 	pipeline_dffe_28;
input 	pipeline_dffe_27;
input 	pipeline_dffe_26;
input 	pipeline_dffe_25;
input 	pipeline_dffe_24;
input 	pipeline_dffe_23;
input 	pipeline_dffe_22;
input 	pipeline_dffe_21;
input 	pipeline_dffe_201;
input 	pipeline_dffe_191;
input 	pipeline_dffe_18;
input 	pipeline_dffe_17;
input 	pipeline_dffe_16;
input 	pipeline_dffe_15;
input 	pipeline_dffe_14;
input 	dxxrv_2;
input 	pipeline_dffe_13;
input 	dxxrv_1;
input 	pipeline_dffe_12;
input 	dxxrv_0;
input 	pipeline_dffe_11;
output 	pipeline_dffe_181;
output 	pipeline_dffe_171;
output 	pipeline_dffe_161;
output 	pipeline_dffe_151;
output 	pipeline_dffe_141;
output 	pipeline_dffe_131;
output 	pipeline_dffe_121;
output 	pipeline_dffe_111;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~82_cout ;
wire \op_1~78_cout ;
wire \op_1~74_cout ;
wire \op_1~70_cout ;
wire \op_1~66 ;
wire \op_1~62 ;
wire \op_1~58 ;
wire \op_1~54 ;
wire \op_1~50 ;
wire \op_1~46 ;
wire \op_1~42 ;
wire \op_1~38 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;


dffeas \pipeline_dffe[19] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \pipeline_dffe[19] .is_wysiwyg = "true";
defparam \pipeline_dffe[19] .power_up = "low";

dffeas \pipeline_dffe[20] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \pipeline_dffe[20] .is_wysiwyg = "true";
defparam \pipeline_dffe[20] .power_up = "low";

dffeas \pipeline_dffe[18] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_181),
	.prn(vcc));
defparam \pipeline_dffe[18] .is_wysiwyg = "true";
defparam \pipeline_dffe[18] .power_up = "low";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_171),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_161),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_151),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_141),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_131),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_121),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_111),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

cyclonev_lcell_comb \op_1~82 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_0),
	.datae(gnd),
	.dataf(!pipeline_dffe_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\op_1~82_cout ),
	.shareout());
defparam \op_1~82 .extended_lut = "off";
defparam \op_1~82 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~82 .shared_arith = "off";

cyclonev_lcell_comb \op_1~78 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_1),
	.datae(gnd),
	.dataf(!pipeline_dffe_12),
	.datag(gnd),
	.cin(\op_1~82_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\op_1~78_cout ),
	.shareout());
defparam \op_1~78 .extended_lut = "off";
defparam \op_1~78 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~78 .shared_arith = "off";

cyclonev_lcell_comb \op_1~74 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_2),
	.datae(gnd),
	.dataf(!pipeline_dffe_13),
	.datag(gnd),
	.cin(\op_1~78_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\op_1~74_cout ),
	.shareout());
defparam \op_1~74 .extended_lut = "off";
defparam \op_1~74 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~74 .shared_arith = "off";

cyclonev_lcell_comb \op_1~70 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_14),
	.datag(gnd),
	.cin(\op_1~74_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\op_1~70_cout ),
	.shareout());
defparam \op_1~70 .extended_lut = "off";
defparam \op_1~70 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~70 .shared_arith = "off";

cyclonev_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_15),
	.datag(gnd),
	.cin(\op_1~70_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

cyclonev_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_16),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

cyclonev_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_17),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

cyclonev_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_18),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

cyclonev_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_191),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_201),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_21),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_22),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_23),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_24),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_25),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_26),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_27),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_28),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_29),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_30),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_31),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

endmodule

module NCO_Lab3_asj_dxx_g (
	dxxrv_3,
	dxxrv_2,
	dxxrv_1,
	dxxrv_0,
	clk,
	reset,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dxxrv_3;
output 	dxxrv_2;
output 	dxxrv_1;
output 	dxxrv_0;
input 	clk;
input 	reset;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lsfr_reg~0_combout ;
wire \lsfr_reg~1_combout ;
wire \lsfr_reg[0]~q ;
wire \lsfr_reg[1]~11_combout ;
wire \lsfr_reg[1]~q ;
wire \lsfr_reg[2]~10_combout ;
wire \lsfr_reg[2]~q ;
wire \lsfr_reg[3]~q ;
wire \lsfr_reg[4]~q ;
wire \lsfr_reg[5]~9_combout ;
wire \lsfr_reg[5]~q ;
wire \lsfr_reg[6]~8_combout ;
wire \lsfr_reg[6]~q ;
wire \lsfr_reg[7]~q ;
wire \lsfr_reg[8]~7_combout ;
wire \lsfr_reg[8]~q ;
wire \lsfr_reg[9]~6_combout ;
wire \lsfr_reg[9]~q ;
wire \lsfr_reg[10]~5_combout ;
wire \lsfr_reg[10]~q ;
wire \lsfr_reg[11]~4_combout ;
wire \lsfr_reg[11]~q ;
wire \lsfr_reg[12]~q ;
wire \lsfr_reg[13]~3_combout ;
wire \lsfr_reg[13]~q ;
wire \lsfr_reg[14]~q ;
wire \lsfr_reg[15]~2_combout ;
wire \lsfr_reg[15]~q ;
wire \Add0~0_combout ;
wire \Add0~1_combout ;
wire \Add0~2_combout ;


dffeas \dxxrv[3] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxrv_3),
	.prn(vcc));
defparam \dxxrv[3] .is_wysiwyg = "true";
defparam \dxxrv[3] .power_up = "low";

dffeas \dxxrv[2] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxrv_2),
	.prn(vcc));
defparam \dxxrv[2] .is_wysiwyg = "true";
defparam \dxxrv[2] .power_up = "low";

dffeas \dxxrv[1] (
	.clk(clk),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxrv_1),
	.prn(vcc));
defparam \dxxrv[1] .is_wysiwyg = "true";
defparam \dxxrv[1] .power_up = "low";

dffeas \dxxrv[0] (
	.clk(clk),
	.d(\lsfr_reg~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dxxrv_0),
	.prn(vcc));
defparam \dxxrv[0] .is_wysiwyg = "true";
defparam \dxxrv[0] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg~0 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~0 .extended_lut = "off";
defparam \lsfr_reg~0 .lut_mask = 64'h6666666666666666;
defparam \lsfr_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \lsfr_reg~1 (
	.dataa(!\lsfr_reg[14]~q ),
	.datab(!\lsfr_reg[3]~q ),
	.datac(!\lsfr_reg~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~1 .extended_lut = "off";
defparam \lsfr_reg~1 .lut_mask = 64'h9696969696969696;
defparam \lsfr_reg~1 .shared_arith = "off";

dffeas \lsfr_reg[0] (
	.clk(clk),
	.d(\lsfr_reg~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[0]~q ),
	.prn(vcc));
defparam \lsfr_reg[0] .is_wysiwyg = "true";
defparam \lsfr_reg[0] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg[1]~11 (
	.dataa(!\lsfr_reg[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg[1]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg[1]~11 .extended_lut = "off";
defparam \lsfr_reg[1]~11 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lsfr_reg[1]~11 .shared_arith = "off";

dffeas \lsfr_reg[1] (
	.clk(clk),
	.d(\lsfr_reg[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[1]~q ),
	.prn(vcc));
defparam \lsfr_reg[1] .is_wysiwyg = "true";
defparam \lsfr_reg[1] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg[2]~10 (
	.dataa(!\lsfr_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg[2]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg[2]~10 .extended_lut = "off";
defparam \lsfr_reg[2]~10 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lsfr_reg[2]~10 .shared_arith = "off";

dffeas \lsfr_reg[2] (
	.clk(clk),
	.d(\lsfr_reg[2]~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[2]~q ),
	.prn(vcc));
defparam \lsfr_reg[2] .is_wysiwyg = "true";
defparam \lsfr_reg[2] .power_up = "low";

dffeas \lsfr_reg[3] (
	.clk(clk),
	.d(\lsfr_reg[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[3]~q ),
	.prn(vcc));
defparam \lsfr_reg[3] .is_wysiwyg = "true";
defparam \lsfr_reg[3] .power_up = "low";

dffeas \lsfr_reg[4] (
	.clk(clk),
	.d(\lsfr_reg[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[4]~q ),
	.prn(vcc));
defparam \lsfr_reg[4] .is_wysiwyg = "true";
defparam \lsfr_reg[4] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg[5]~9 (
	.dataa(!\lsfr_reg[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg[5]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg[5]~9 .extended_lut = "off";
defparam \lsfr_reg[5]~9 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lsfr_reg[5]~9 .shared_arith = "off";

dffeas \lsfr_reg[5] (
	.clk(clk),
	.d(\lsfr_reg[5]~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[5]~q ),
	.prn(vcc));
defparam \lsfr_reg[5] .is_wysiwyg = "true";
defparam \lsfr_reg[5] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg[6]~8 (
	.dataa(!\lsfr_reg[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg[6]~8 .extended_lut = "off";
defparam \lsfr_reg[6]~8 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lsfr_reg[6]~8 .shared_arith = "off";

dffeas \lsfr_reg[6] (
	.clk(clk),
	.d(\lsfr_reg[6]~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[6]~q ),
	.prn(vcc));
defparam \lsfr_reg[6] .is_wysiwyg = "true";
defparam \lsfr_reg[6] .power_up = "low";

dffeas \lsfr_reg[7] (
	.clk(clk),
	.d(\lsfr_reg[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[7]~q ),
	.prn(vcc));
defparam \lsfr_reg[7] .is_wysiwyg = "true";
defparam \lsfr_reg[7] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg[8]~7 (
	.dataa(!\lsfr_reg[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg[8]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg[8]~7 .extended_lut = "off";
defparam \lsfr_reg[8]~7 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lsfr_reg[8]~7 .shared_arith = "off";

dffeas \lsfr_reg[8] (
	.clk(clk),
	.d(\lsfr_reg[8]~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[8]~q ),
	.prn(vcc));
defparam \lsfr_reg[8] .is_wysiwyg = "true";
defparam \lsfr_reg[8] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg[9]~6 (
	.dataa(!\lsfr_reg[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg[9]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg[9]~6 .extended_lut = "off";
defparam \lsfr_reg[9]~6 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lsfr_reg[9]~6 .shared_arith = "off";

dffeas \lsfr_reg[9] (
	.clk(clk),
	.d(\lsfr_reg[9]~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[9]~q ),
	.prn(vcc));
defparam \lsfr_reg[9] .is_wysiwyg = "true";
defparam \lsfr_reg[9] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg[10]~5 (
	.dataa(!\lsfr_reg[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg[10]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg[10]~5 .extended_lut = "off";
defparam \lsfr_reg[10]~5 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lsfr_reg[10]~5 .shared_arith = "off";

dffeas \lsfr_reg[10] (
	.clk(clk),
	.d(\lsfr_reg[10]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[10]~q ),
	.prn(vcc));
defparam \lsfr_reg[10] .is_wysiwyg = "true";
defparam \lsfr_reg[10] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg[11]~4 (
	.dataa(!\lsfr_reg[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg[11]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg[11]~4 .extended_lut = "off";
defparam \lsfr_reg[11]~4 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lsfr_reg[11]~4 .shared_arith = "off";

dffeas \lsfr_reg[11] (
	.clk(clk),
	.d(\lsfr_reg[11]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[11]~q ),
	.prn(vcc));
defparam \lsfr_reg[11] .is_wysiwyg = "true";
defparam \lsfr_reg[11] .power_up = "low";

dffeas \lsfr_reg[12] (
	.clk(clk),
	.d(\lsfr_reg[11]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[12]~q ),
	.prn(vcc));
defparam \lsfr_reg[12] .is_wysiwyg = "true";
defparam \lsfr_reg[12] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg[13]~3 (
	.dataa(!\lsfr_reg[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg[13]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg[13]~3 .extended_lut = "off";
defparam \lsfr_reg[13]~3 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lsfr_reg[13]~3 .shared_arith = "off";

dffeas \lsfr_reg[13] (
	.clk(clk),
	.d(\lsfr_reg[13]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[13]~q ),
	.prn(vcc));
defparam \lsfr_reg[13] .is_wysiwyg = "true";
defparam \lsfr_reg[13] .power_up = "low";

dffeas \lsfr_reg[14] (
	.clk(clk),
	.d(\lsfr_reg[13]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[14]~q ),
	.prn(vcc));
defparam \lsfr_reg[14] .is_wysiwyg = "true";
defparam \lsfr_reg[14] .power_up = "low";

cyclonev_lcell_comb \lsfr_reg[15]~2 (
	.dataa(!\lsfr_reg[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg[15]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg[15]~2 .extended_lut = "off";
defparam \lsfr_reg[15]~2 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \lsfr_reg[15]~2 .shared_arith = "off";

dffeas \lsfr_reg[15] (
	.clk(clk),
	.d(\lsfr_reg[15]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\lsfr_reg[15]~q ),
	.prn(vcc));
defparam \lsfr_reg[15] .is_wysiwyg = "true";
defparam \lsfr_reg[15] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[14]~q ),
	.datac(!\lsfr_reg[13]~q ),
	.datad(!\lsfr_reg[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \Add0~0 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[14]~q ),
	.datac(!\lsfr_reg[13]~q ),
	.datad(!\lsfr_reg[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h6996699669966996;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~2 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[13]~q ),
	.datac(!\lsfr_reg[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~2 .extended_lut = "off";
defparam \Add0~2 .lut_mask = 64'h9696969696969696;
defparam \Add0~2 .shared_arith = "off";

endmodule

module NCO_Lab3_asj_nco_isdr (
	data_ready1,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	data_ready1;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lpm_counter_component|auto_generated|counter_reg_bit[1]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[0]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[4]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[3]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[2]~q ;
wire \always0~0_combout ;
wire \data_ready~0_combout ;


NCO_Lab3_lpm_counter_1 lpm_counter_component(
	.counter_reg_bit_1(\lpm_counter_component|auto_generated|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\lpm_counter_component|auto_generated|counter_reg_bit[0]~q ),
	.counter_reg_bit_4(\lpm_counter_component|auto_generated|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\lpm_counter_component|auto_generated|counter_reg_bit[3]~q ),
	.counter_reg_bit_2(\lpm_counter_component|auto_generated|counter_reg_bit[2]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas data_ready(
	.clk(clk),
	.d(\data_ready~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_ready1),
	.prn(vcc));
defparam data_ready.is_wysiwyg = "true";
defparam data_ready.power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!clken),
	.datab(!\lpm_counter_component|auto_generated|counter_reg_bit[4]~q ),
	.datac(!\lpm_counter_component|auto_generated|counter_reg_bit[3]~q ),
	.datad(!\lpm_counter_component|auto_generated|counter_reg_bit[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \data_ready~0 (
	.dataa(!data_ready1),
	.datab(!\lpm_counter_component|auto_generated|counter_reg_bit[1]~q ),
	.datac(!\lpm_counter_component|auto_generated|counter_reg_bit[0]~q ),
	.datad(!\always0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_ready~0 .extended_lut = "off";
defparam \data_ready~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \data_ready~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_counter_1 (
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_cntr_bki auto_generated(
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.counter_reg_bit_2(counter_reg_bit_2),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_cntr_bki (
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_4,
	counter_reg_bit_3,
	counter_reg_bit_2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
output 	counter_reg_bit_2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita3~sumout ;
wire \counter_comb_bita2~sumout ;


dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

cyclonev_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

cyclonev_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

endmodule

module NCO_Lab3_cord_2c (
	cordic_x_res_2c_0,
	cordic_y_res_2c_0,
	cordic_y_res_d_1,
	cordic_x_res_d_1,
	cordic_y_res_2c_1,
	cordic_x_res_2c_1,
	cordic_y_res_d_2,
	cordic_x_res_d_2,
	cordic_y_res_2c_2,
	cordic_x_res_2c_2,
	cordic_y_res_d_3,
	cordic_x_res_d_3,
	cordic_y_res_2c_3,
	cordic_x_res_2c_3,
	cordic_y_res_d_4,
	cordic_x_res_d_4,
	cordic_y_res_2c_4,
	cordic_x_res_2c_4,
	cordic_y_res_d_5,
	cordic_x_res_d_5,
	cordic_y_res_2c_5,
	cordic_x_res_2c_5,
	cordic_y_res_d_6,
	cordic_x_res_d_6,
	cordic_y_res_2c_6,
	cordic_x_res_2c_6,
	cordic_y_res_d_7,
	cordic_x_res_d_7,
	cordic_y_res_2c_7,
	cordic_x_res_2c_7,
	cordic_y_res_d_8,
	cordic_x_res_d_8,
	cordic_y_res_2c_8,
	cordic_x_res_2c_8,
	cordic_y_res_d_9,
	cordic_x_res_d_9,
	cordic_y_res_2c_9,
	cordic_x_res_2c_9,
	cordic_y_res_d_10,
	cordic_x_res_d_10,
	cordic_y_res_2c_10,
	cordic_x_res_2c_10,
	cordic_y_res_d_11,
	cordic_x_res_d_11,
	cordic_y_res_2c_11,
	cordic_x_res_2c_11,
	dffe1,
	pipeline_dffe_0,
	pipeline_dffe_1,
	dffe2,
	pipeline_dffe_2,
	dffe3,
	pipeline_dffe_3,
	dffe4,
	pipeline_dffe_4,
	dffe5,
	pipeline_dffe_5,
	dffe6,
	pipeline_dffe_6,
	dffe7,
	pipeline_dffe_7,
	dffe8,
	pipeline_dffe_8,
	dffe9,
	pipeline_dffe_9,
	dffe10,
	pipeline_dffe_10,
	dffe11,
	pipeline_dffe_11,
	dffe12,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	cordic_x_res_2c_0;
output 	cordic_y_res_2c_0;
output 	cordic_y_res_d_1;
output 	cordic_x_res_d_1;
output 	cordic_y_res_2c_1;
output 	cordic_x_res_2c_1;
output 	cordic_y_res_d_2;
output 	cordic_x_res_d_2;
output 	cordic_y_res_2c_2;
output 	cordic_x_res_2c_2;
output 	cordic_y_res_d_3;
output 	cordic_x_res_d_3;
output 	cordic_y_res_2c_3;
output 	cordic_x_res_2c_3;
output 	cordic_y_res_d_4;
output 	cordic_x_res_d_4;
output 	cordic_y_res_2c_4;
output 	cordic_x_res_2c_4;
output 	cordic_y_res_d_5;
output 	cordic_x_res_d_5;
output 	cordic_y_res_2c_5;
output 	cordic_x_res_2c_5;
output 	cordic_y_res_d_6;
output 	cordic_x_res_d_6;
output 	cordic_y_res_2c_6;
output 	cordic_x_res_2c_6;
output 	cordic_y_res_d_7;
output 	cordic_x_res_d_7;
output 	cordic_y_res_2c_7;
output 	cordic_x_res_2c_7;
output 	cordic_y_res_d_8;
output 	cordic_x_res_d_8;
output 	cordic_y_res_2c_8;
output 	cordic_x_res_2c_8;
output 	cordic_y_res_d_9;
output 	cordic_x_res_d_9;
output 	cordic_y_res_2c_9;
output 	cordic_x_res_2c_9;
output 	cordic_y_res_d_10;
output 	cordic_x_res_d_10;
output 	cordic_y_res_2c_10;
output 	cordic_x_res_2c_10;
output 	cordic_y_res_d_11;
output 	cordic_x_res_d_11;
output 	cordic_y_res_2c_11;
output 	cordic_x_res_2c_11;
input 	dffe1;
input 	pipeline_dffe_0;
input 	pipeline_dffe_1;
input 	dffe2;
input 	pipeline_dffe_2;
input 	dffe3;
input 	pipeline_dffe_3;
input 	dffe4;
input 	pipeline_dffe_4;
input 	dffe5;
input 	pipeline_dffe_5;
input 	dffe6;
input 	pipeline_dffe_6;
input 	dffe7;
input 	pipeline_dffe_7;
input 	dffe8;
input 	pipeline_dffe_8;
input 	dffe9;
input 	pipeline_dffe_9;
input 	dffe10;
input 	pipeline_dffe_10;
input 	dffe11;
input 	pipeline_dffe_11;
input 	dffe12;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add1~1_sumout ;
wire \Add0~1_sumout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add1~22 ;
wire \Add1~25_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add1~26 ;
wire \Add1~29_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add1~30 ;
wire \Add1~33_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add1~34 ;
wire \Add1~37_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add1~38 ;
wire \Add1~41_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;


dffeas \cordic_x_res_2c[0] (
	.clk(clk),
	.d(dffe1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_0),
	.prn(vcc));
defparam \cordic_x_res_2c[0] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[0] .power_up = "low";

dffeas \cordic_y_res_2c[0] (
	.clk(clk),
	.d(pipeline_dffe_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_0),
	.prn(vcc));
defparam \cordic_y_res_2c[0] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[0] .power_up = "low";

dffeas \cordic_y_res_d[1] (
	.clk(clk),
	.d(pipeline_dffe_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_1),
	.prn(vcc));
defparam \cordic_y_res_d[1] .is_wysiwyg = "true";
defparam \cordic_y_res_d[1] .power_up = "low";

dffeas \cordic_x_res_d[1] (
	.clk(clk),
	.d(dffe2),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_1),
	.prn(vcc));
defparam \cordic_x_res_d[1] .is_wysiwyg = "true";
defparam \cordic_x_res_d[1] .power_up = "low";

dffeas \cordic_y_res_2c[1] (
	.clk(clk),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_1),
	.prn(vcc));
defparam \cordic_y_res_2c[1] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[1] .power_up = "low";

dffeas \cordic_x_res_2c[1] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_1),
	.prn(vcc));
defparam \cordic_x_res_2c[1] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[1] .power_up = "low";

dffeas \cordic_y_res_d[2] (
	.clk(clk),
	.d(pipeline_dffe_2),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_2),
	.prn(vcc));
defparam \cordic_y_res_d[2] .is_wysiwyg = "true";
defparam \cordic_y_res_d[2] .power_up = "low";

dffeas \cordic_x_res_d[2] (
	.clk(clk),
	.d(dffe3),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_2),
	.prn(vcc));
defparam \cordic_x_res_d[2] .is_wysiwyg = "true";
defparam \cordic_x_res_d[2] .power_up = "low";

dffeas \cordic_y_res_2c[2] (
	.clk(clk),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_2),
	.prn(vcc));
defparam \cordic_y_res_2c[2] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[2] .power_up = "low";

dffeas \cordic_x_res_2c[2] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_2),
	.prn(vcc));
defparam \cordic_x_res_2c[2] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[2] .power_up = "low";

dffeas \cordic_y_res_d[3] (
	.clk(clk),
	.d(pipeline_dffe_3),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_3),
	.prn(vcc));
defparam \cordic_y_res_d[3] .is_wysiwyg = "true";
defparam \cordic_y_res_d[3] .power_up = "low";

dffeas \cordic_x_res_d[3] (
	.clk(clk),
	.d(dffe4),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_3),
	.prn(vcc));
defparam \cordic_x_res_d[3] .is_wysiwyg = "true";
defparam \cordic_x_res_d[3] .power_up = "low";

dffeas \cordic_y_res_2c[3] (
	.clk(clk),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_3),
	.prn(vcc));
defparam \cordic_y_res_2c[3] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[3] .power_up = "low";

dffeas \cordic_x_res_2c[3] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_3),
	.prn(vcc));
defparam \cordic_x_res_2c[3] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[3] .power_up = "low";

dffeas \cordic_y_res_d[4] (
	.clk(clk),
	.d(pipeline_dffe_4),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_4),
	.prn(vcc));
defparam \cordic_y_res_d[4] .is_wysiwyg = "true";
defparam \cordic_y_res_d[4] .power_up = "low";

dffeas \cordic_x_res_d[4] (
	.clk(clk),
	.d(dffe5),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_4),
	.prn(vcc));
defparam \cordic_x_res_d[4] .is_wysiwyg = "true";
defparam \cordic_x_res_d[4] .power_up = "low";

dffeas \cordic_y_res_2c[4] (
	.clk(clk),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_4),
	.prn(vcc));
defparam \cordic_y_res_2c[4] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[4] .power_up = "low";

dffeas \cordic_x_res_2c[4] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_4),
	.prn(vcc));
defparam \cordic_x_res_2c[4] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[4] .power_up = "low";

dffeas \cordic_y_res_d[5] (
	.clk(clk),
	.d(pipeline_dffe_5),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_5),
	.prn(vcc));
defparam \cordic_y_res_d[5] .is_wysiwyg = "true";
defparam \cordic_y_res_d[5] .power_up = "low";

dffeas \cordic_x_res_d[5] (
	.clk(clk),
	.d(dffe6),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_5),
	.prn(vcc));
defparam \cordic_x_res_d[5] .is_wysiwyg = "true";
defparam \cordic_x_res_d[5] .power_up = "low";

dffeas \cordic_y_res_2c[5] (
	.clk(clk),
	.d(\Add1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_5),
	.prn(vcc));
defparam \cordic_y_res_2c[5] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[5] .power_up = "low";

dffeas \cordic_x_res_2c[5] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_5),
	.prn(vcc));
defparam \cordic_x_res_2c[5] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[5] .power_up = "low";

dffeas \cordic_y_res_d[6] (
	.clk(clk),
	.d(pipeline_dffe_6),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_6),
	.prn(vcc));
defparam \cordic_y_res_d[6] .is_wysiwyg = "true";
defparam \cordic_y_res_d[6] .power_up = "low";

dffeas \cordic_x_res_d[6] (
	.clk(clk),
	.d(dffe7),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_6),
	.prn(vcc));
defparam \cordic_x_res_d[6] .is_wysiwyg = "true";
defparam \cordic_x_res_d[6] .power_up = "low";

dffeas \cordic_y_res_2c[6] (
	.clk(clk),
	.d(\Add1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_6),
	.prn(vcc));
defparam \cordic_y_res_2c[6] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[6] .power_up = "low";

dffeas \cordic_x_res_2c[6] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_6),
	.prn(vcc));
defparam \cordic_x_res_2c[6] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[6] .power_up = "low";

dffeas \cordic_y_res_d[7] (
	.clk(clk),
	.d(pipeline_dffe_7),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_7),
	.prn(vcc));
defparam \cordic_y_res_d[7] .is_wysiwyg = "true";
defparam \cordic_y_res_d[7] .power_up = "low";

dffeas \cordic_x_res_d[7] (
	.clk(clk),
	.d(dffe8),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_7),
	.prn(vcc));
defparam \cordic_x_res_d[7] .is_wysiwyg = "true";
defparam \cordic_x_res_d[7] .power_up = "low";

dffeas \cordic_y_res_2c[7] (
	.clk(clk),
	.d(\Add1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_7),
	.prn(vcc));
defparam \cordic_y_res_2c[7] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[7] .power_up = "low";

dffeas \cordic_x_res_2c[7] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_7),
	.prn(vcc));
defparam \cordic_x_res_2c[7] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[7] .power_up = "low";

dffeas \cordic_y_res_d[8] (
	.clk(clk),
	.d(pipeline_dffe_8),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_8),
	.prn(vcc));
defparam \cordic_y_res_d[8] .is_wysiwyg = "true";
defparam \cordic_y_res_d[8] .power_up = "low";

dffeas \cordic_x_res_d[8] (
	.clk(clk),
	.d(dffe9),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_8),
	.prn(vcc));
defparam \cordic_x_res_d[8] .is_wysiwyg = "true";
defparam \cordic_x_res_d[8] .power_up = "low";

dffeas \cordic_y_res_2c[8] (
	.clk(clk),
	.d(\Add1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_8),
	.prn(vcc));
defparam \cordic_y_res_2c[8] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[8] .power_up = "low";

dffeas \cordic_x_res_2c[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_8),
	.prn(vcc));
defparam \cordic_x_res_2c[8] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[8] .power_up = "low";

dffeas \cordic_y_res_d[9] (
	.clk(clk),
	.d(pipeline_dffe_9),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_9),
	.prn(vcc));
defparam \cordic_y_res_d[9] .is_wysiwyg = "true";
defparam \cordic_y_res_d[9] .power_up = "low";

dffeas \cordic_x_res_d[9] (
	.clk(clk),
	.d(dffe10),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_9),
	.prn(vcc));
defparam \cordic_x_res_d[9] .is_wysiwyg = "true";
defparam \cordic_x_res_d[9] .power_up = "low";

dffeas \cordic_y_res_2c[9] (
	.clk(clk),
	.d(\Add1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_9),
	.prn(vcc));
defparam \cordic_y_res_2c[9] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[9] .power_up = "low";

dffeas \cordic_x_res_2c[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_9),
	.prn(vcc));
defparam \cordic_x_res_2c[9] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[9] .power_up = "low";

dffeas \cordic_y_res_d[10] (
	.clk(clk),
	.d(pipeline_dffe_10),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_10),
	.prn(vcc));
defparam \cordic_y_res_d[10] .is_wysiwyg = "true";
defparam \cordic_y_res_d[10] .power_up = "low";

dffeas \cordic_x_res_d[10] (
	.clk(clk),
	.d(dffe11),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_10),
	.prn(vcc));
defparam \cordic_x_res_d[10] .is_wysiwyg = "true";
defparam \cordic_x_res_d[10] .power_up = "low";

dffeas \cordic_y_res_2c[10] (
	.clk(clk),
	.d(\Add1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_10),
	.prn(vcc));
defparam \cordic_y_res_2c[10] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[10] .power_up = "low";

dffeas \cordic_x_res_2c[10] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_10),
	.prn(vcc));
defparam \cordic_x_res_2c[10] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[10] .power_up = "low";

dffeas \cordic_y_res_d[11] (
	.clk(clk),
	.d(pipeline_dffe_11),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_d_11),
	.prn(vcc));
defparam \cordic_y_res_d[11] .is_wysiwyg = "true";
defparam \cordic_y_res_d[11] .power_up = "low";

dffeas \cordic_x_res_d[11] (
	.clk(clk),
	.d(dffe12),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_d_11),
	.prn(vcc));
defparam \cordic_x_res_d[11] .is_wysiwyg = "true";
defparam \cordic_x_res_d[11] .power_up = "low";

dffeas \cordic_y_res_2c[11] (
	.clk(clk),
	.d(\Add1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_y_res_2c_11),
	.prn(vcc));
defparam \cordic_y_res_2c[11] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[11] .power_up = "low";

dffeas \cordic_x_res_2c[11] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cordic_x_res_2c_11),
	.prn(vcc));
defparam \cordic_x_res_2c[11] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[11] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_0),
	.datae(gnd),
	.dataf(!pipeline_dffe_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000FF0000FF00;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe2),
	.datae(gnd),
	.dataf(!dffe1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000000000FF00;
defparam \Add1~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000000000FF00;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000000000FF00;
defparam \Add1~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000000000FF00;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000000000FF00;
defparam \Add1~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000000000FF00;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h000000000000FF00;
defparam \Add1~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000000000FF00;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h000000000000FF00;
defparam \Add1~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000000000FF00;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000000000FF00;
defparam \Add1~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h000000000000FF00;
defparam \Add1~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000000000FF00;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout());
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h000000000000FF00;
defparam \Add1~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000000000FF00;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~37_sumout ),
	.cout(\Add1~38 ),
	.shareout());
defparam \Add1~37 .extended_lut = "off";
defparam \Add1~37 .lut_mask = 64'h000000000000FF00;
defparam \Add1~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000000000FF00;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~41_sumout ),
	.cout(),
	.shareout());
defparam \Add1~41 .extended_lut = "off";
defparam \Add1~41 .lut_mask = 64'h000000000000FF00;
defparam \Add1~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000000000FF00;
defparam \Add0~41 .shared_arith = "off";

endmodule

module NCO_Lab3_cord_fs (
	cor1x_10,
	corx_10,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	cor1x_10;
input 	corx_10;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \cor1x[10] (
	.clk(clk),
	.d(corx_10),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(cor1x_10),
	.prn(vcc));
defparam \cor1x[10] .is_wysiwyg = "true";
defparam \cor1x[10] .power_up = "low";

endmodule

module NCO_Lab3_cord_init (
	corx_10,
	corz_14,
	dxxpdo_18,
	corz_13,
	dxxpdo_17,
	corz_12,
	dxxpdo_16,
	corz_11,
	dxxpdo_15,
	corz_10,
	dxxpdo_14,
	corz_9,
	dxxpdo_13,
	corz_8,
	dxxpdo_12,
	corz_7,
	dxxpdo_11,
	corz_6,
	dxxpdo_10,
	corz_5,
	dxxpdo_9,
	corz_4,
	dxxpdo_8,
	corz_3,
	dxxpdo_7,
	corz_2,
	dxxpdo_6,
	corz_1,
	dxxpdo_5,
	corz_0,
	dxxpdo_4,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	corx_10;
output 	corz_14;
input 	dxxpdo_18;
output 	corz_13;
input 	dxxpdo_17;
output 	corz_12;
input 	dxxpdo_16;
output 	corz_11;
input 	dxxpdo_15;
output 	corz_10;
input 	dxxpdo_14;
output 	corz_9;
input 	dxxpdo_13;
output 	corz_8;
input 	dxxpdo_12;
output 	corz_7;
input 	dxxpdo_11;
output 	corz_6;
input 	dxxpdo_10;
output 	corz_5;
input 	dxxpdo_9;
output 	corz_4;
input 	dxxpdo_8;
output 	corz_3;
input 	dxxpdo_7;
output 	corz_2;
input 	dxxpdo_6;
output 	corz_1;
input 	dxxpdo_5;
output 	corz_0;
input 	dxxpdo_4;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \corx[10] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corx_10),
	.prn(vcc));
defparam \corx[10] .is_wysiwyg = "true";
defparam \corx[10] .power_up = "low";

dffeas \corz[14] (
	.clk(clk),
	.d(dxxpdo_18),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_14),
	.prn(vcc));
defparam \corz[14] .is_wysiwyg = "true";
defparam \corz[14] .power_up = "low";

dffeas \corz[13] (
	.clk(clk),
	.d(dxxpdo_17),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_13),
	.prn(vcc));
defparam \corz[13] .is_wysiwyg = "true";
defparam \corz[13] .power_up = "low";

dffeas \corz[12] (
	.clk(clk),
	.d(dxxpdo_16),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_12),
	.prn(vcc));
defparam \corz[12] .is_wysiwyg = "true";
defparam \corz[12] .power_up = "low";

dffeas \corz[11] (
	.clk(clk),
	.d(dxxpdo_15),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_11),
	.prn(vcc));
defparam \corz[11] .is_wysiwyg = "true";
defparam \corz[11] .power_up = "low";

dffeas \corz[10] (
	.clk(clk),
	.d(dxxpdo_14),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_10),
	.prn(vcc));
defparam \corz[10] .is_wysiwyg = "true";
defparam \corz[10] .power_up = "low";

dffeas \corz[9] (
	.clk(clk),
	.d(dxxpdo_13),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_9),
	.prn(vcc));
defparam \corz[9] .is_wysiwyg = "true";
defparam \corz[9] .power_up = "low";

dffeas \corz[8] (
	.clk(clk),
	.d(dxxpdo_12),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_8),
	.prn(vcc));
defparam \corz[8] .is_wysiwyg = "true";
defparam \corz[8] .power_up = "low";

dffeas \corz[7] (
	.clk(clk),
	.d(dxxpdo_11),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_7),
	.prn(vcc));
defparam \corz[7] .is_wysiwyg = "true";
defparam \corz[7] .power_up = "low";

dffeas \corz[6] (
	.clk(clk),
	.d(dxxpdo_10),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_6),
	.prn(vcc));
defparam \corz[6] .is_wysiwyg = "true";
defparam \corz[6] .power_up = "low";

dffeas \corz[5] (
	.clk(clk),
	.d(dxxpdo_9),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_5),
	.prn(vcc));
defparam \corz[5] .is_wysiwyg = "true";
defparam \corz[5] .power_up = "low";

dffeas \corz[4] (
	.clk(clk),
	.d(dxxpdo_8),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_4),
	.prn(vcc));
defparam \corz[4] .is_wysiwyg = "true";
defparam \corz[4] .power_up = "low";

dffeas \corz[3] (
	.clk(clk),
	.d(dxxpdo_7),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_3),
	.prn(vcc));
defparam \corz[3] .is_wysiwyg = "true";
defparam \corz[3] .power_up = "low";

dffeas \corz[2] (
	.clk(clk),
	.d(dxxpdo_6),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_2),
	.prn(vcc));
defparam \corz[2] .is_wysiwyg = "true";
defparam \corz[2] .power_up = "low";

dffeas \corz[1] (
	.clk(clk),
	.d(dxxpdo_5),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_1),
	.prn(vcc));
defparam \corz[1] .is_wysiwyg = "true";
defparam \corz[1] .power_up = "low";

dffeas \corz[0] (
	.clk(clk),
	.d(dxxpdo_4),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(corz_0),
	.prn(vcc));
defparam \corz[0] .is_wysiwyg = "true";
defparam \corz[0] .power_up = "low";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm (
	pipeline_dffe_11,
	pipeline_dffe_10,
	dffe16,
	pipeline_dffe_9,
	pipeline_dffe_111,
	dffe12,
	pipeline_dffe_8,
	pipeline_dffe_7,
	dffe11,
	pipeline_dffe_101,
	pipeline_dffe_6,
	dffe10,
	pipeline_dffe_91,
	pipeline_dffe_4,
	pipeline_dffe_5,
	dffe9,
	pipeline_dffe_81,
	dffe8,
	pipeline_dffe_71,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	dffe7,
	pipeline_dffe_61,
	dffe6,
	pipeline_dffe_51,
	pipeline_dffe_31,
	pipeline_dffe_41,
	dffe5,
	dffe4,
	pipeline_dffe_01,
	pipeline_dffe_12,
	pipeline_dffe_21,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	dffe16;
output 	pipeline_dffe_9;
input 	pipeline_dffe_111;
input 	dffe12;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
input 	dffe11;
input 	pipeline_dffe_101;
output 	pipeline_dffe_6;
input 	dffe10;
input 	pipeline_dffe_91;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
input 	dffe9;
input 	pipeline_dffe_81;
input 	dffe8;
input 	pipeline_dffe_71;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
input 	dffe7;
input 	pipeline_dffe_61;
input 	dffe6;
input 	pipeline_dffe_51;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	dffe5;
input 	dffe4;
input 	pipeline_dffe_01;
input 	pipeline_dffe_12;
input 	pipeline_dffe_21;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \xordvalue~1_combout ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \xordvalue~2_combout ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \xordvalue[0]~q ;
wire \a[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;


NCO_Lab3_lpm_add_sub_3 u0(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_10(\a[10]~q ),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_9(\a[9]~q ),
	.pipeline_dffe_7(pipeline_dffe_7),
	.a_8(\a[8]~q ),
	.pipeline_dffe_6(pipeline_dffe_6),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_0(\a[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!dffe8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

cyclonev_lcell_comb \xordvalue~5 (
	.dataa(!dffe7),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~6 (
	.dataa(!dffe4),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~7 (
	.dataa(!dffe5),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~8 (
	.dataa(!dffe6),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_3 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	pipeline_dffe_9,
	a_10,
	pipeline_dffe_8,
	a_9,
	pipeline_dffe_7,
	a_8,
	pipeline_dffe_6,
	a_7,
	xordvalue_7,
	pipeline_dffe_4,
	pipeline_dffe_5,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	a_4,
	xordvalue_4,
	a_3,
	xordvalue_3,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_9;
input 	a_10;
output 	pipeline_dffe_8;
input 	a_9;
output 	pipeline_dffe_7;
input 	a_8;
output 	pipeline_dffe_6;
input 	a_7;
input 	xordvalue_7;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
input 	a_4;
input 	xordvalue_4;
input 	a_3;
input 	xordvalue_3;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_10(a_10),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_9(a_9),
	.pipeline_dffe_7(pipeline_dffe_7),
	.a_8(a_8),
	.pipeline_dffe_6(pipeline_dffe_6),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.xordvalue_0(xordvalue_0),
	.a_0(a_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h (
	pipeline_dffe_11,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	pipeline_dffe_9,
	a_10,
	pipeline_dffe_8,
	a_9,
	pipeline_dffe_7,
	a_8,
	pipeline_dffe_6,
	a_7,
	xordvalue_7,
	pipeline_dffe_4,
	pipeline_dffe_5,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	a_4,
	xordvalue_4,
	a_3,
	xordvalue_3,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_9;
input 	a_10;
output 	pipeline_dffe_8;
input 	a_9;
output 	pipeline_dffe_7;
input 	a_8;
output 	pipeline_dffe_6;
input 	a_7;
input 	xordvalue_7;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
input 	a_4;
input 	xordvalue_4;
input 	a_3;
input 	xordvalue_3;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~29_sumout ;
wire \op_1~25_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~33_sumout ;


dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm_1 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	dffe16,
	dffe12,
	pipeline_dffe_9,
	pipeline_dffe_111,
	pipeline_dffe_8,
	pipeline_dffe_101,
	pipeline_dffe_7,
	dffe11,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_91,
	dffe10,
	pipeline_dffe_81,
	dffe9,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_71,
	dffe8,
	pipeline_dffe_61,
	dffe7,
	pipeline_dffe_41,
	pipeline_dffe_51,
	dffe6,
	dffe5,
	pipeline_dffe_01,
	pipeline_dffe_12,
	pipeline_dffe_21,
	pipeline_dffe_31,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	dffe16;
input 	dffe12;
output 	pipeline_dffe_9;
input 	pipeline_dffe_111;
output 	pipeline_dffe_8;
input 	pipeline_dffe_101;
output 	pipeline_dffe_7;
input 	dffe11;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
input 	pipeline_dffe_91;
input 	dffe10;
input 	pipeline_dffe_81;
input 	dffe9;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
input 	pipeline_dffe_71;
input 	dffe8;
input 	pipeline_dffe_61;
input 	dffe7;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	dffe6;
input 	dffe5;
input 	pipeline_dffe_01;
input 	pipeline_dffe_12;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \xordvalue[0]~q ;
wire \a[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;


NCO_Lab3_lpm_add_sub_4 u0(
	.pipeline_dffe_11(pipeline_dffe_11),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_10(\a[10]~q ),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_9(\a[9]~q ),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_8(\a[8]~q ),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_0(\a[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!dffe9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!dffe5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!dffe6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!dffe7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!dffe8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_4 (
	pipeline_dffe_11,
	a_11,
	xordvalue_10,
	pipeline_dffe_10,
	a_10,
	pipeline_dffe_9,
	a_9,
	pipeline_dffe_8,
	a_8,
	pipeline_dffe_7,
	pipeline_dffe_5,
	pipeline_dffe_6,
	a_7,
	a_6,
	xordvalue_6,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_10;
input 	a_10;
output 	pipeline_dffe_9;
input 	a_9;
output 	pipeline_dffe_8;
input 	a_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
input 	a_7;
input 	a_6;
input 	xordvalue_6;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h_1 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_10(a_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_9(a_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_8(a_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.a_7(a_7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.xordvalue_0(xordvalue_0),
	.a_0(a_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h_1 (
	pipeline_dffe_11,
	a_11,
	xordvalue_10,
	pipeline_dffe_10,
	a_10,
	pipeline_dffe_9,
	a_9,
	pipeline_dffe_8,
	a_8,
	pipeline_dffe_7,
	pipeline_dffe_5,
	pipeline_dffe_6,
	a_7,
	a_6,
	xordvalue_6,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_10;
input 	a_10;
output 	pipeline_dffe_9;
input 	a_9;
output 	pipeline_dffe_8;
input 	a_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
input 	a_7;
input 	a_6;
input 	xordvalue_6;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~25_sumout ;
wire \op_1~21_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~29_sumout ;


dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm_2 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	dffe16,
	pipeline_dffe_9,
	pipeline_dffe_111,
	dffe12,
	pipeline_dffe_8,
	pipeline_dffe_6,
	pipeline_dffe_7,
	dffe11,
	pipeline_dffe_101,
	dffe10,
	pipeline_dffe_91,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	dffe9,
	pipeline_dffe_81,
	dffe8,
	pipeline_dffe_71,
	pipeline_dffe_51,
	pipeline_dffe_61,
	dffe7,
	dffe6,
	pipeline_dffe_01,
	pipeline_dffe_12,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	dffe16;
output 	pipeline_dffe_9;
input 	pipeline_dffe_111;
input 	dffe12;
output 	pipeline_dffe_8;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	dffe11;
input 	pipeline_dffe_101;
input 	dffe10;
input 	pipeline_dffe_91;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
input 	dffe9;
input 	pipeline_dffe_81;
input 	dffe8;
input 	pipeline_dffe_71;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	dffe7;
input 	dffe6;
input 	pipeline_dffe_01;
input 	pipeline_dffe_12;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \xordvalue[0]~q ;
wire \a[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;


NCO_Lab3_lpm_add_sub_5 u0(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_10(\a[10]~q ),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_9(\a[9]~q ),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_0(\a[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe6),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe7),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!dffe8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~5 (
	.dataa(!dffe9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~6 (
	.dataa(!dffe10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_5 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	pipeline_dffe_9,
	a_10,
	pipeline_dffe_8,
	a_9,
	pipeline_dffe_6,
	pipeline_dffe_7,
	a_8,
	a_7,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	a_6,
	a_5,
	xordvalue_5,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_9;
input 	a_10;
output 	pipeline_dffe_8;
input 	a_9;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	a_8;
input 	a_7;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
input 	a_6;
input 	a_5;
input 	xordvalue_5;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h_2 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_10(a_10),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_9(a_9),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.a_8(a_8),
	.a_7(a_7),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.a_6(a_6),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.xordvalue_0(xordvalue_0),
	.a_0(a_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h_2 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	pipeline_dffe_9,
	a_10,
	pipeline_dffe_8,
	a_9,
	pipeline_dffe_6,
	pipeline_dffe_7,
	a_8,
	a_7,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	a_6,
	a_5,
	xordvalue_5,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_9;
input 	a_10;
output 	pipeline_dffe_8;
input 	a_9;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	a_8;
input 	a_7;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
input 	a_6;
input 	a_5;
input 	xordvalue_5;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~21_sumout ;
wire \op_1~17_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~25_sumout ;


dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm_3 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	dffe16,
	dffe12,
	pipeline_dffe_9,
	pipeline_dffe_111,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_101,
	dffe11,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_91,
	dffe10,
	pipeline_dffe_81,
	dffe9,
	pipeline_dffe_61,
	pipeline_dffe_71,
	dffe8,
	dffe7,
	pipeline_dffe_01,
	pipeline_dffe_12,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	dffe16;
input 	dffe12;
output 	pipeline_dffe_9;
input 	pipeline_dffe_111;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	pipeline_dffe_101;
input 	dffe11;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
input 	pipeline_dffe_91;
input 	dffe10;
input 	pipeline_dffe_81;
input 	dffe9;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	dffe8;
input 	dffe7;
input 	pipeline_dffe_01;
input 	pipeline_dffe_12;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \xordvalue[0]~q ;
wire \a[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;


NCO_Lab3_lpm_add_sub_6 u0(
	.pipeline_dffe_11(pipeline_dffe_11),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_10(\a[10]~q ),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_0(\a[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!dffe9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!dffe10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!dffe11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_6 (
	pipeline_dffe_11,
	a_11,
	xordvalue_10,
	pipeline_dffe_10,
	a_10,
	pipeline_dffe_9,
	pipeline_dffe_7,
	pipeline_dffe_8,
	a_9,
	a_8,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	a_7,
	a_6,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_10;
input 	a_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	a_9;
input 	a_8;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
input 	a_7;
input 	a_6;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h_3 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_10(a_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_9(a_9),
	.a_8(a_8),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.a_7(a_7),
	.a_6(a_6),
	.xordvalue_0(xordvalue_0),
	.a_0(a_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h_3 (
	pipeline_dffe_11,
	a_11,
	xordvalue_10,
	pipeline_dffe_10,
	a_10,
	pipeline_dffe_9,
	pipeline_dffe_7,
	pipeline_dffe_8,
	a_9,
	a_8,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	a_7,
	a_6,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_10;
input 	a_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	a_9;
input 	a_8;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
input 	a_7;
input 	a_6;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~26 ;
wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~17_sumout ;
wire \op_1~13_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~21_sumout ;


dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm_4 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_8,
	pipeline_dffe_9,
	dffe16,
	pipeline_dffe_111,
	dffe12,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	dffe11,
	pipeline_dffe_101,
	dffe10,
	pipeline_dffe_91,
	pipeline_dffe_71,
	pipeline_dffe_81,
	dffe9,
	dffe8,
	pipeline_dffe_01,
	pipeline_dffe_12,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	dffe16;
input 	pipeline_dffe_111;
input 	dffe12;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	dffe11;
input 	pipeline_dffe_101;
input 	dffe10;
input 	pipeline_dffe_91;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	dffe9;
input 	dffe8;
input 	pipeline_dffe_01;
input 	pipeline_dffe_12;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \xordvalue[0]~q ;
wire \a[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;


NCO_Lab3_lpm_add_sub_7 u0(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_0(\a[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!dffe11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_7 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	pipeline_dffe_8,
	pipeline_dffe_9,
	a_10,
	a_9,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	a_8,
	a_7,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	a_5,
	a_6,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	a_10;
input 	a_9;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	a_8;
input 	a_7;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h_4 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_10(a_10),
	.a_9(a_9),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.a_8(a_8),
	.a_7(a_7),
	.xordvalue_0(xordvalue_0),
	.a_0(a_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h_4 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	pipeline_dffe_8,
	pipeline_dffe_9,
	a_10,
	a_9,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	a_8,
	a_7,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	a_5,
	a_6,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	a_10;
input 	a_9;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	a_8;
input 	a_7;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~22 ;
wire \op_1~26 ;
wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~13_sumout ;
wire \op_1~9_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~17_sumout ;


dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm_5 (
	pipeline_dffe_11,
	pipeline_dffe_9,
	pipeline_dffe_10,
	dffe16,
	dffe12,
	pipeline_dffe_111,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_101,
	dffe11,
	pipeline_dffe_81,
	pipeline_dffe_91,
	dffe10,
	dffe9,
	pipeline_dffe_01,
	pipeline_dffe_12,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
input 	dffe16;
input 	dffe12;
input 	pipeline_dffe_111;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	pipeline_dffe_101;
input 	dffe11;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	dffe10;
input 	dffe9;
input 	pipeline_dffe_01;
input 	pipeline_dffe_12;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \xordvalue[0]~q ;
wire \a[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;


NCO_Lab3_lpm_add_sub_8 u0(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_10(\a[10]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_0(\a[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!dffe11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_8 (
	pipeline_dffe_11,
	pipeline_dffe_9,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	a_10,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	a_9,
	a_8,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
input 	a_10;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	a_9;
input 	a_8;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h_5 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.a_10(a_10),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_9(a_9),
	.a_8(a_8),
	.xordvalue_0(xordvalue_0),
	.a_0(a_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h_5 (
	pipeline_dffe_11,
	pipeline_dffe_9,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	a_10,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	a_9,
	a_8,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
input 	a_10;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	a_9;
input 	a_8;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~18 ;
wire \op_1~22 ;
wire \op_1~26 ;
wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~9_sumout ;
wire \op_1~5_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~13_sumout ;


dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm_6 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	dffe16,
	pipeline_dffe_111,
	dffe12,
	pipeline_dffe_91,
	pipeline_dffe_101,
	dffe11,
	dffe10,
	pipeline_dffe_01,
	pipeline_dffe_12,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	dffe16;
input 	pipeline_dffe_111;
input 	dffe12;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	dffe11;
input 	dffe10;
input 	pipeline_dffe_01;
input 	pipeline_dffe_12;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \a[10]~q ;
wire \xordvalue~0_combout ;
wire \a[9]~q ;
wire \xordvalue[0]~q ;
wire \a[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;


NCO_Lab3_lpm_add_sub_9 u0(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_0(\a[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_9 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	a_10,
	a_9,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	a_10;
input 	a_9;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h_6 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_10(a_10),
	.a_9(a_9),
	.xordvalue_0(xordvalue_0),
	.a_0(a_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h_6 (
	pipeline_dffe_11,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	a_10,
	a_9,
	xordvalue_0,
	a_0,
	a_1,
	xordvalue_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	a_10;
input 	a_9;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~14 ;
wire \op_1~18 ;
wire \op_1~22 ;
wire \op_1~26 ;
wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~9_sumout ;


dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm_7 (
	pipeline_dffe_11,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	dffe16,
	dffe12,
	pipeline_dffe_111,
	pipeline_dffe_101,
	dffe11,
	pipeline_dffe_01,
	pipeline_dffe_12,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
input 	dffe16;
input 	dffe12;
input 	pipeline_dffe_111;
input 	pipeline_dffe_101;
input 	dffe11;
input 	pipeline_dffe_01;
input 	pipeline_dffe_12;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \xordvalue[0]~q ;
wire \a[0]~q ;
wire \a[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \xordvalue~1_combout ;


NCO_Lab3_lpm_add_sub_10 u0(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_0(\a[0]~q ),
	.a_1(\a[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_10 (
	pipeline_dffe_11,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	a_10,
	xordvalue_0,
	a_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
input 	a_10;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h_7 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.a_10(a_10),
	.xordvalue_0(xordvalue_0),
	.a_0(a_0),
	.a_1(a_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h_7 (
	pipeline_dffe_11,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	a_11,
	xordvalue_10,
	a_10,
	xordvalue_0,
	a_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
input 	a_11;
input 	xordvalue_10;
input 	a_10;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~10 ;
wire \op_1~14 ;
wire \op_1~18 ;
wire \op_1~22 ;
wire \op_1~26 ;
wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~5_sumout ;


dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm_8 (
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	dffe16,
	pipeline_dffe_111,
	dffe12,
	pipeline_dffe_01,
	pipeline_dffe_12,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	dffe16;
input 	pipeline_dffe_111;
input 	dffe12;
input 	pipeline_dffe_01;
input 	pipeline_dffe_12;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \xordvalue[0]~q ;
wire \a[0]~q ;
wire \a[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \xordvalue~0_combout ;


NCO_Lab3_lpm_add_sub_11 u0(
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_0(\a[0]~q ),
	.a_1(\a[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_11 (
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	xordvalue_0,
	a_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h_8 auto_generated(
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.xordvalue_0(xordvalue_0),
	.a_0(a_0),
	.a_1(a_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h_8 (
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	xordvalue_0,
	a_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	xordvalue_0;
input 	a_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~30 ;
wire \op_1~33_sumout ;
wire \op_1~34 ;
wire \op_1~37_sumout ;
wire \op_1~38 ;
wire \op_1~41_sumout ;
wire \op_1~42 ;
wire \op_1~45_sumout ;


dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_1),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_2),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_3),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_4),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_5),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_6),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_7),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_8),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_9),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_10),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_11),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm_9 (
	pipeline_dffe_11,
	a_0,
	xordvalue_2,
	pipeline_dffe_10,
	dffe16,
	cor1x_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	a_0;
output 	xordvalue_2;
output 	pipeline_dffe_10;
input 	dffe16;
input 	cor1x_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[10]~q ;
wire \xordvalue~0_combout ;


NCO_Lab3_lpm_add_sub_12 u0(
	.pipeline_dffe_11(pipeline_dffe_11),
	.a_0(a_0),
	.xordvalue_2(xordvalue_2),
	.a_10(\a[10]~q ),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[10] (
	.clk(clk),
	.d(cor1x_10),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(dffe16),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(a_0),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(xordvalue_2),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!cor1x_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_12 (
	pipeline_dffe_11,
	a_0,
	xordvalue_2,
	a_10,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
input 	a_0;
input 	xordvalue_2;
input 	a_10;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h_9 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.a_0(a_0),
	.xordvalue_2(xordvalue_2),
	.a_10(a_10),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h_9 (
	pipeline_dffe_11,
	a_0,
	xordvalue_2,
	a_10,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
input 	a_0;
input 	xordvalue_2;
input 	a_10;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~0_combout ;
wire \op_1~1_combout ;
wire \op_1~2_combout ;
wire \op_1~3_combout ;
wire \op_1~4_combout ;
wire \op_1~5_combout ;
wire \op_1~6_combout ;
wire \op_1~7_combout ;
wire \op_1~8_combout ;


dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

cyclonev_lcell_comb \op_1~0 (
	.dataa(!a_0),
	.datab(!xordvalue_2),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~0 .extended_lut = "off";
defparam \op_1~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \op_1~0 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(!a_0),
	.datab(!xordvalue_2),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h9696969696969696;
defparam \op_1~1 .shared_arith = "off";

cyclonev_lcell_comb \op_1~2 (
	.dataa(!a_0),
	.datab(!xordvalue_2),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~2 .extended_lut = "off";
defparam \op_1~2 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \op_1~2 .shared_arith = "off";

cyclonev_lcell_comb \op_1~3 (
	.dataa(!a_0),
	.datab(!xordvalue_2),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~3 .extended_lut = "off";
defparam \op_1~3 .lut_mask = 64'h9696969696969696;
defparam \op_1~3 .shared_arith = "off";

cyclonev_lcell_comb \op_1~4 (
	.dataa(!a_0),
	.datab(!xordvalue_2),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~4 .extended_lut = "off";
defparam \op_1~4 .lut_mask = 64'h9696969696969696;
defparam \op_1~4 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(!a_0),
	.datab(!xordvalue_2),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~6 (
	.dataa(!a_0),
	.datab(!xordvalue_2),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~6 .extended_lut = "off";
defparam \op_1~6 .lut_mask = 64'h9696969696969696;
defparam \op_1~6 .shared_arith = "off";

cyclonev_lcell_comb \op_1~7 (
	.dataa(!a_0),
	.datab(!xordvalue_2),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~7 .extended_lut = "off";
defparam \op_1~7 .lut_mask = 64'h9696969696969696;
defparam \op_1~7 .shared_arith = "off";

cyclonev_lcell_comb \op_1~8 (
	.dataa(!a_0),
	.datab(!xordvalue_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~8 .extended_lut = "off";
defparam \op_1~8 .lut_mask = 64'h6666666666666666;
defparam \op_1~8 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_axor_1p_lpm_10 (
	pipeline_dffe_11,
	a_0,
	pipeline_dffe_10,
	dffe16,
	pipeline_dffe_111,
	dffe12,
	pipeline_dffe_9,
	pipeline_dffe_101,
	pipeline_dffe_8,
	pipeline_dffe_91,
	pipeline_dffe_7,
	dffe11,
	pipeline_dffe_81,
	pipeline_dffe_6,
	dffe10,
	pipeline_dffe_71,
	pipeline_dffe_5,
	dffe9,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_61,
	dffe8,
	pipeline_dffe_51,
	dffe7,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_41,
	dffe6,
	pipeline_dffe_31,
	dffe5,
	pipeline_dffe_21,
	dffe4,
	dffe3,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
output 	a_0;
output 	pipeline_dffe_10;
input 	dffe16;
input 	pipeline_dffe_111;
input 	dffe12;
output 	pipeline_dffe_9;
input 	pipeline_dffe_101;
output 	pipeline_dffe_8;
input 	pipeline_dffe_91;
output 	pipeline_dffe_7;
input 	dffe11;
input 	pipeline_dffe_81;
output 	pipeline_dffe_6;
input 	dffe10;
input 	pipeline_dffe_71;
output 	pipeline_dffe_5;
input 	dffe9;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
input 	pipeline_dffe_61;
input 	dffe8;
input 	pipeline_dffe_51;
input 	dffe7;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
input 	pipeline_dffe_41;
input 	dffe6;
input 	pipeline_dffe_31;
input 	dffe5;
input 	pipeline_dffe_21;
input 	dffe4;
input 	dffe3;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \xordvalue~1_combout ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \xordvalue~2_combout ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \xordvalue~3_combout ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \xordvalue~4_combout ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \xordvalue[0]~q ;
wire \xordvalue[1]~q ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;


NCO_Lab3_lpm_add_sub_13 u0(
	.pipeline_dffe_11(pipeline_dffe_11),
	.a_0(a_0),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_10(\a[10]~q ),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_9(\a[9]~q ),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.pipeline_dffe_7(pipeline_dffe_7),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.pipeline_dffe_6(pipeline_dffe_6),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[11] (
	.clk(clk),
	.d(pipeline_dffe_111),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(pipeline_dffe_101),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(pipeline_dffe_91),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(pipeline_dffe_81),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

dffeas \a[7] (
	.clk(clk),
	.d(pipeline_dffe_71),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

dffeas \a[6] (
	.clk(clk),
	.d(pipeline_dffe_61),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!dffe9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

dffeas \a[5] (
	.clk(clk),
	.d(pipeline_dffe_51),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!dffe8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

dffeas \a[4] (
	.clk(clk),
	.d(pipeline_dffe_41),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(pipeline_dffe_31),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

cyclonev_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!dffe7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!dffe6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

dffeas \a[2] (
	.clk(clk),
	.d(pipeline_dffe_21),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

cyclonev_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!dffe5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!dffe3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~9 (
	.dataa(!dffe16),
	.datab(!dffe4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

dffeas \a[0] (
	.clk(clk),
	.d(dffe16),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(a_0),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

endmodule

module NCO_Lab3_lpm_add_sub_13 (
	pipeline_dffe_11,
	a_0,
	a_11,
	xordvalue_10,
	pipeline_dffe_10,
	a_10,
	pipeline_dffe_9,
	a_9,
	pipeline_dffe_8,
	a_8,
	xordvalue_8,
	pipeline_dffe_7,
	a_7,
	xordvalue_7,
	pipeline_dffe_6,
	a_6,
	xordvalue_6,
	pipeline_dffe_5,
	pipeline_dffe_3,
	pipeline_dffe_4,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	a_3,
	xordvalue_3,
	a_2,
	xordvalue_2,
	xordvalue_0,
	xordvalue_1,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
input 	a_0;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_10;
input 	a_10;
output 	pipeline_dffe_9;
input 	a_9;
output 	pipeline_dffe_8;
input 	a_8;
input 	xordvalue_8;
output 	pipeline_dffe_7;
input 	a_7;
input 	xordvalue_7;
output 	pipeline_dffe_6;
input 	a_6;
input 	xordvalue_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
input 	a_3;
input 	xordvalue_3;
input 	a_2;
input 	xordvalue_2;
input 	xordvalue_0;
input 	xordvalue_1;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_o0h_10 auto_generated(
	.pipeline_dffe_11(pipeline_dffe_11),
	.a_0(a_0),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.pipeline_dffe_10(pipeline_dffe_10),
	.a_10(a_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.a_9(a_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.xordvalue_0(xordvalue_0),
	.xordvalue_1(xordvalue_1),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_o0h_10 (
	pipeline_dffe_11,
	a_0,
	a_11,
	xordvalue_10,
	pipeline_dffe_10,
	a_10,
	pipeline_dffe_9,
	a_9,
	pipeline_dffe_8,
	a_8,
	xordvalue_8,
	pipeline_dffe_7,
	a_7,
	xordvalue_7,
	pipeline_dffe_6,
	a_6,
	xordvalue_6,
	pipeline_dffe_5,
	pipeline_dffe_3,
	pipeline_dffe_4,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	a_3,
	xordvalue_3,
	a_2,
	xordvalue_2,
	xordvalue_0,
	xordvalue_1,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_11;
input 	a_0;
input 	a_11;
input 	xordvalue_10;
output 	pipeline_dffe_10;
input 	a_10;
output 	pipeline_dffe_9;
input 	a_9;
output 	pipeline_dffe_8;
input 	a_8;
input 	xordvalue_8;
output 	pipeline_dffe_7;
input 	a_7;
input 	xordvalue_7;
output 	pipeline_dffe_6;
input 	a_6;
input 	xordvalue_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
input 	a_3;
input 	xordvalue_3;
input 	a_2;
input 	xordvalue_2;
input 	xordvalue_0;
input 	xordvalue_1;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~38 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~33_sumout ;
wire \op_1~29_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~37_sumout ;


dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

cyclonev_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

cyclonev_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h00000000000000FF;
defparam \op_1~45 .shared_arith = "off";

cyclonev_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

cyclonev_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

cyclonev_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

cyclonev_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

cyclonev_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

cyclonev_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

cyclonev_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

cyclonev_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

cyclonev_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

cyclonev_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm (
	dffe12,
	dffe11,
	dffe16,
	pipeline_dffe_11,
	dffe10,
	dffe121,
	dffe9,
	dffe111,
	dffe8,
	pipeline_dffe_10,
	dffe101,
	dffe7,
	pipeline_dffe_9,
	dffe91,
	dffe6,
	pipeline_dffe_8,
	dffe5,
	dffe1,
	dffe81,
	pipeline_dffe_7,
	dffe2,
	dffe3,
	dffe4,
	dffe71,
	pipeline_dffe_6,
	dffe61,
	pipeline_dffe_5,
	pipeline_dffe_3,
	pipeline_dffe_4,
	dffe51,
	dffe41,
	dffe13,
	dffe21,
	dffe31,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
input 	dffe16;
input 	pipeline_dffe_11;
output 	dffe10;
input 	dffe121;
output 	dffe9;
input 	dffe111;
output 	dffe8;
input 	pipeline_dffe_10;
input 	dffe101;
output 	dffe7;
input 	pipeline_dffe_9;
input 	dffe91;
output 	dffe6;
input 	pipeline_dffe_8;
output 	dffe5;
output 	dffe1;
input 	dffe81;
input 	pipeline_dffe_7;
output 	dffe2;
output 	dffe3;
output 	dffe4;
input 	dffe71;
input 	pipeline_dffe_6;
input 	dffe61;
input 	pipeline_dffe_5;
input 	pipeline_dffe_3;
input 	pipeline_dffe_4;
input 	dffe51;
input 	dffe41;
input 	dffe13;
input 	dffe21;
input 	dffe31;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \xordvalue~1_combout ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \xordvalue~2_combout ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \xordvalue~3_combout ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \xordvalue~4_combout ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;


NCO_Lab3_lpm_add_sub_14 u0(
	.dffe12(dffe12),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe11(dffe11),
	.a_10(\a[10]~q ),
	.dffe10(dffe10),
	.a_9(\a[9]~q ),
	.dffe9(dffe9),
	.a_8(\a[8]~q ),
	.dffe8(dffe8),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.dffe7(dffe7),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe1(dffe1),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe13),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

cyclonev_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_14 (
	dffe12,
	a_11,
	xordvalue_10,
	dffe11,
	a_10,
	dffe10,
	a_9,
	dffe9,
	a_8,
	dffe8,
	a_7,
	xordvalue_7,
	dffe7,
	a_6,
	xordvalue_6,
	dffe6,
	dffe5,
	dffe1,
	a_5,
	xordvalue_5,
	dffe2,
	dffe3,
	dffe4,
	a_4,
	xordvalue_4,
	a_0,
	xordvalue_0,
	a_3,
	xordvalue_3,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
input 	a_11;
input 	xordvalue_10;
output 	dffe11;
input 	a_10;
output 	dffe10;
input 	a_9;
output 	dffe9;
input 	a_8;
output 	dffe8;
input 	a_7;
input 	xordvalue_7;
output 	dffe7;
input 	a_6;
input 	xordvalue_6;
output 	dffe6;
output 	dffe5;
output 	dffe1;
input 	a_5;
input 	xordvalue_5;
output 	dffe2;
output 	dffe3;
output 	dffe4;
input 	a_4;
input 	xordvalue_4;
input 	a_0;
input 	xordvalue_0;
input 	a_3;
input 	xordvalue_3;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg auto_generated(
	.dffe121(dffe12),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.dffe111(dffe11),
	.a_10(a_10),
	.dffe101(dffe10),
	.a_9(a_9),
	.dffe91(dffe9),
	.a_8(a_8),
	.dffe81(dffe8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.dffe71(dffe7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe13(dffe1),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg (
	dffe121,
	a_11,
	xordvalue_10,
	dffe111,
	a_10,
	dffe101,
	a_9,
	dffe91,
	a_8,
	dffe81,
	a_7,
	xordvalue_7,
	dffe71,
	a_6,
	xordvalue_6,
	dffe61,
	dffe51,
	dffe13,
	a_5,
	xordvalue_5,
	dffe21,
	dffe31,
	dffe41,
	a_4,
	xordvalue_4,
	a_0,
	xordvalue_0,
	a_3,
	xordvalue_3,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe121;
input 	a_11;
input 	xordvalue_10;
output 	dffe111;
input 	a_10;
output 	dffe101;
input 	a_9;
output 	dffe91;
input 	a_8;
output 	dffe81;
input 	a_7;
input 	xordvalue_7;
output 	dffe71;
input 	a_6;
input 	xordvalue_6;
output 	dffe61;
output 	dffe51;
output 	dffe13;
input 	a_5;
input 	xordvalue_5;
output 	dffe21;
output 	dffe31;
output 	dffe41;
input 	a_4;
input 	xordvalue_4;
input 	a_0;
input 	xordvalue_0;
input 	a_3;
input 	xordvalue_3;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;


dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm_1 (
	dffe12,
	dffe11,
	dffe16,
	dffe10,
	dffe121,
	pipeline_dffe_11,
	dffe9,
	dffe8,
	pipeline_dffe_10,
	dffe111,
	dffe7,
	pipeline_dffe_9,
	dffe101,
	dffe6,
	dffe1,
	pipeline_dffe_8,
	dffe91,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	pipeline_dffe_7,
	dffe81,
	pipeline_dffe_6,
	dffe71,
	pipeline_dffe_4,
	pipeline_dffe_5,
	dffe61,
	dffe51,
	dffe13,
	dffe21,
	dffe31,
	dffe41,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
input 	dffe16;
output 	dffe10;
input 	dffe121;
input 	pipeline_dffe_11;
output 	dffe9;
output 	dffe8;
input 	pipeline_dffe_10;
input 	dffe111;
output 	dffe7;
input 	pipeline_dffe_9;
input 	dffe101;
output 	dffe6;
output 	dffe1;
input 	pipeline_dffe_8;
input 	dffe91;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
input 	pipeline_dffe_7;
input 	dffe81;
input 	pipeline_dffe_6;
input 	dffe71;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	dffe61;
input 	dffe51;
input 	dffe13;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \xordvalue~1_combout ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \xordvalue~2_combout ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;


NCO_Lab3_lpm_add_sub_15 u0(
	.dffe12(dffe12),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.dffe6(dffe6),
	.dffe1(dffe1),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe13),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!pipeline_dffe_9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!pipeline_dffe_4),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!pipeline_dffe_8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~5 (
	.dataa(!pipeline_dffe_5),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~6 (
	.dataa(!pipeline_dffe_6),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~7 (
	.dataa(!pipeline_dffe_7),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_15 (
	dffe12,
	dffe11,
	a_11,
	xordvalue_10,
	dffe10,
	a_10,
	dffe9,
	a_9,
	dffe8,
	a_8,
	dffe7,
	a_7,
	dffe6,
	dffe1,
	a_6,
	xordvalue_6,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	a_5,
	xordvalue_5,
	a_0,
	xordvalue_0,
	a_4,
	xordvalue_4,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
input 	a_11;
input 	xordvalue_10;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
input 	a_8;
output 	dffe7;
input 	a_7;
output 	dffe6;
output 	dffe1;
input 	a_6;
input 	xordvalue_6;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
input 	a_5;
input 	xordvalue_5;
input 	a_0;
input 	xordvalue_0;
input 	a_4;
input 	xordvalue_4;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg_1 auto_generated(
	.dffe121(dffe12),
	.dffe111(dffe11),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.a_8(a_8),
	.dffe71(dffe7),
	.a_7(a_7),
	.dffe61(dffe6),
	.dffe13(dffe1),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg_1 (
	dffe121,
	dffe111,
	a_11,
	xordvalue_10,
	dffe101,
	a_10,
	dffe91,
	a_9,
	dffe81,
	a_8,
	dffe71,
	a_7,
	dffe61,
	dffe13,
	a_6,
	xordvalue_6,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	a_5,
	xordvalue_5,
	a_0,
	xordvalue_0,
	a_4,
	xordvalue_4,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe121;
output 	dffe111;
input 	a_11;
input 	xordvalue_10;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
input 	a_8;
output 	dffe71;
input 	a_7;
output 	dffe61;
output 	dffe13;
input 	a_6;
input 	xordvalue_6;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
input 	a_5;
input 	xordvalue_5;
input 	a_0;
input 	xordvalue_0;
input 	a_4;
input 	xordvalue_4;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;


dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm_2 (
	dffe12,
	dffe11,
	dffe16,
	pipeline_dffe_11,
	dffe10,
	dffe121,
	dffe9,
	dffe111,
	dffe8,
	pipeline_dffe_10,
	dffe7,
	dffe1,
	dffe101,
	pipeline_dffe_9,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe91,
	pipeline_dffe_8,
	dffe81,
	pipeline_dffe_7,
	pipeline_dffe_5,
	pipeline_dffe_6,
	dffe71,
	dffe61,
	dffe13,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
input 	dffe16;
input 	pipeline_dffe_11;
output 	dffe10;
input 	dffe121;
output 	dffe9;
input 	dffe111;
output 	dffe8;
input 	pipeline_dffe_10;
output 	dffe7;
output 	dffe1;
input 	dffe101;
input 	pipeline_dffe_9;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
input 	dffe91;
input 	pipeline_dffe_8;
input 	dffe81;
input 	pipeline_dffe_7;
input 	pipeline_dffe_5;
input 	pipeline_dffe_6;
input 	dffe71;
input 	dffe61;
input 	dffe13;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;


NCO_Lab3_lpm_add_sub_16 u0(
	.dffe12(dffe12),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe11(dffe11),
	.a_10(\a[10]~q ),
	.dffe10(dffe10),
	.a_9(\a[9]~q ),
	.dffe9(dffe9),
	.a_8(\a[8]~q ),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe1(dffe1),
	.a_7(\a[7]~q ),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe13),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_16 (
	dffe12,
	a_11,
	xordvalue_10,
	dffe11,
	a_10,
	dffe10,
	a_9,
	dffe9,
	a_8,
	dffe8,
	dffe7,
	dffe1,
	a_7,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	a_6,
	a_0,
	xordvalue_0,
	a_5,
	xordvalue_5,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
input 	a_11;
input 	xordvalue_10;
output 	dffe11;
input 	a_10;
output 	dffe10;
input 	a_9;
output 	dffe9;
input 	a_8;
output 	dffe8;
output 	dffe7;
output 	dffe1;
input 	a_7;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
input 	a_6;
input 	a_0;
input 	xordvalue_0;
input 	a_5;
input 	xordvalue_5;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg_2 auto_generated(
	.dffe121(dffe12),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.dffe111(dffe11),
	.a_10(a_10),
	.dffe101(dffe10),
	.a_9(a_9),
	.dffe91(dffe9),
	.a_8(a_8),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe13(dffe1),
	.a_7(a_7),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.a_6(a_6),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg_2 (
	dffe121,
	a_11,
	xordvalue_10,
	dffe111,
	a_10,
	dffe101,
	a_9,
	dffe91,
	a_8,
	dffe81,
	dffe71,
	dffe13,
	a_7,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	a_6,
	a_0,
	xordvalue_0,
	a_5,
	xordvalue_5,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe121;
input 	a_11;
input 	xordvalue_10;
output 	dffe111;
input 	a_10;
output 	dffe101;
input 	a_9;
output 	dffe91;
input 	a_8;
output 	dffe81;
output 	dffe71;
output 	dffe13;
input 	a_7;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
input 	a_6;
input 	a_0;
input 	xordvalue_0;
input 	a_5;
input 	xordvalue_5;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;


dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm_3 (
	dffe12,
	dffe11,
	dffe16,
	dffe10,
	dffe121,
	pipeline_dffe_11,
	dffe9,
	dffe8,
	dffe1,
	pipeline_dffe_10,
	dffe111,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	pipeline_dffe_9,
	dffe101,
	pipeline_dffe_8,
	dffe91,
	pipeline_dffe_6,
	pipeline_dffe_7,
	dffe81,
	dffe71,
	dffe13,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
input 	dffe16;
output 	dffe10;
input 	dffe121;
input 	pipeline_dffe_11;
output 	dffe9;
output 	dffe8;
output 	dffe1;
input 	pipeline_dffe_10;
input 	dffe111;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
input 	pipeline_dffe_9;
input 	dffe101;
input 	pipeline_dffe_8;
input 	dffe91;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	dffe81;
input 	dffe71;
input 	dffe13;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[6]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;


NCO_Lab3_lpm_add_sub_17 u0(
	.dffe12(dffe12),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.dffe1(dffe1),
	.a_8(\a[8]~q ),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_6(\a[6]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe13),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_6),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!pipeline_dffe_7),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!pipeline_dffe_8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!pipeline_dffe_9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~5 (
	.dataa(!pipeline_dffe_10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_17 (
	dffe12,
	dffe11,
	a_11,
	xordvalue_10,
	dffe10,
	a_10,
	dffe9,
	a_9,
	dffe8,
	dffe1,
	a_8,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	a_7,
	a_0,
	xordvalue_0,
	a_6,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
input 	a_11;
input 	xordvalue_10;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
output 	dffe1;
input 	a_8;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
input 	a_7;
input 	a_0;
input 	xordvalue_0;
input 	a_6;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg_3 auto_generated(
	.dffe121(dffe12),
	.dffe111(dffe11),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.dffe13(dffe1),
	.a_8(a_8),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.a_7(a_7),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_6(a_6),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg_3 (
	dffe121,
	dffe111,
	a_11,
	xordvalue_10,
	dffe101,
	a_10,
	dffe91,
	a_9,
	dffe81,
	dffe13,
	a_8,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	a_7,
	a_0,
	xordvalue_0,
	a_6,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe121;
output 	dffe111;
input 	a_11;
input 	xordvalue_10;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
output 	dffe13;
input 	a_8;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
input 	a_7;
input 	a_0;
input 	xordvalue_0;
input 	a_6;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;


dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm_4 (
	dffe12,
	dffe11,
	dffe16,
	pipeline_dffe_11,
	dffe10,
	dffe121,
	dffe9,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe111,
	pipeline_dffe_10,
	dffe101,
	pipeline_dffe_9,
	pipeline_dffe_7,
	pipeline_dffe_8,
	dffe91,
	dffe81,
	dffe13,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
input 	dffe16;
input 	pipeline_dffe_11;
output 	dffe10;
input 	dffe121;
output 	dffe9;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
input 	dffe111;
input 	pipeline_dffe_10;
input 	dffe101;
input 	pipeline_dffe_9;
input 	pipeline_dffe_7;
input 	pipeline_dffe_8;
input 	dffe91;
input 	dffe81;
input 	dffe13;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[7]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;


NCO_Lab3_lpm_add_sub_18 u0(
	.dffe12(dffe12),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe11(dffe11),
	.a_10(\a[10]~q ),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe1(dffe1),
	.a_9(\a[9]~q ),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_7(\a[7]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe13),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_18 (
	dffe12,
	a_11,
	xordvalue_10,
	dffe11,
	a_10,
	dffe10,
	dffe9,
	dffe1,
	a_9,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	a_8,
	a_0,
	xordvalue_0,
	a_7,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	a_5,
	a_6,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
input 	a_11;
input 	xordvalue_10;
output 	dffe11;
input 	a_10;
output 	dffe10;
output 	dffe9;
output 	dffe1;
input 	a_9;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
input 	a_8;
input 	a_0;
input 	xordvalue_0;
input 	a_7;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg_4 auto_generated(
	.dffe121(dffe12),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.dffe111(dffe11),
	.a_10(a_10),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe13(dffe1),
	.a_9(a_9),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.a_8(a_8),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_7(a_7),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg_4 (
	dffe121,
	a_11,
	xordvalue_10,
	dffe111,
	a_10,
	dffe101,
	dffe91,
	dffe13,
	a_9,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	a_8,
	a_0,
	xordvalue_0,
	a_7,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	a_5,
	a_6,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe121;
input 	a_11;
input 	xordvalue_10;
output 	dffe111;
input 	a_10;
output 	dffe101;
output 	dffe91;
output 	dffe13;
input 	a_9;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
input 	a_8;
input 	a_0;
input 	xordvalue_0;
input 	a_7;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;


dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm_5 (
	dffe12,
	dffe11,
	dffe10,
	dffe1,
	dffe16,
	dffe121,
	pipeline_dffe_11,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	pipeline_dffe_10,
	dffe111,
	pipeline_dffe_8,
	pipeline_dffe_9,
	dffe101,
	dffe91,
	dffe13,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe1;
input 	dffe16;
input 	dffe121;
input 	pipeline_dffe_11;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
input 	pipeline_dffe_10;
input 	dffe111;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	dffe101;
input 	dffe91;
input 	dffe13;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[8]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;


NCO_Lab3_lpm_add_sub_19 u0(
	.dffe12(dffe12),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe10(dffe10),
	.dffe1(dffe1),
	.a_10(\a[10]~q ),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_8(\a[8]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe13),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!pipeline_dffe_9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!pipeline_dffe_10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_19 (
	dffe12,
	dffe11,
	a_11,
	xordvalue_10,
	dffe10,
	dffe1,
	a_10,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	a_9,
	a_0,
	xordvalue_0,
	a_8,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
input 	a_11;
input 	xordvalue_10;
output 	dffe10;
output 	dffe1;
input 	a_10;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
input 	a_9;
input 	a_0;
input 	xordvalue_0;
input 	a_8;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg_5 auto_generated(
	.dffe121(dffe12),
	.dffe111(dffe11),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.dffe101(dffe10),
	.dffe13(dffe1),
	.a_10(a_10),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.a_9(a_9),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_8(a_8),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg_5 (
	dffe121,
	dffe111,
	a_11,
	xordvalue_10,
	dffe101,
	dffe13,
	a_10,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	a_9,
	a_0,
	xordvalue_0,
	a_8,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe121;
output 	dffe111;
input 	a_11;
input 	xordvalue_10;
output 	dffe101;
output 	dffe13;
input 	a_10;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
input 	a_9;
input 	a_0;
input 	xordvalue_0;
input 	a_8;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;


dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm_6 (
	dffe12,
	dffe11,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe16,
	pipeline_dffe_11,
	dffe121,
	pipeline_dffe_9,
	pipeline_dffe_10,
	dffe111,
	dffe101,
	dffe13,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
input 	dffe16;
input 	pipeline_dffe_11;
input 	dffe121;
input 	pipeline_dffe_9;
input 	pipeline_dffe_10;
input 	dffe111;
input 	dffe101;
input 	dffe13;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[9]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;


NCO_Lab3_lpm_add_sub_20 u0(
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe1(dffe1),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_9(\a[9]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe13),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_20 (
	dffe12,
	dffe11,
	dffe1,
	a_11,
	xordvalue_10,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	a_10,
	a_0,
	xordvalue_0,
	a_9,
	a_1,
	xordvalue_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
output 	dffe1;
input 	a_11;
input 	xordvalue_10;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
input 	a_10;
input 	a_0;
input 	xordvalue_0;
input 	a_9;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg_6 auto_generated(
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe13(dffe1),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.a_10(a_10),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_9(a_9),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg_6 (
	dffe121,
	dffe111,
	dffe13,
	a_11,
	xordvalue_10,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	a_10,
	a_0,
	xordvalue_0,
	a_9,
	a_1,
	xordvalue_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe121;
output 	dffe111;
output 	dffe13;
input 	a_11;
input 	xordvalue_10;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
input 	a_10;
input 	a_0;
input 	xordvalue_0;
input 	a_9;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;


dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm_7 (
	dffe12,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe16,
	dffe121,
	pipeline_dffe_11,
	pipeline_dffe_10,
	dffe111,
	dffe13,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
input 	dffe16;
input 	dffe121;
input 	pipeline_dffe_11;
input 	pipeline_dffe_10;
input 	dffe111;
input 	dffe13;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	dffe101;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \xordvalue~1_combout ;


NCO_Lab3_lpm_add_sub_21 u0(
	.dffe12(dffe12),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_10(\a[10]~q ),
	.a_1(\a[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe13),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_21 (
	dffe12,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	a_11,
	xordvalue_10,
	a_0,
	xordvalue_0,
	a_10,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
input 	a_11;
input 	xordvalue_10;
input 	a_0;
input 	xordvalue_0;
input 	a_10;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg_7 auto_generated(
	.dffe121(dffe12),
	.dffe13(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_10(a_10),
	.a_1(a_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg_7 (
	dffe121,
	dffe13,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	a_11,
	xordvalue_10,
	a_0,
	xordvalue_0,
	a_10,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe121;
output 	dffe13;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
output 	dffe111;
input 	a_11;
input 	xordvalue_10;
input 	a_0;
input 	xordvalue_0;
input 	a_10;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[10]~sumout ;


dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm_8 (
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe16,
	pipeline_dffe_11,
	dffe121,
	dffe13,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
input 	dffe16;
input 	pipeline_dffe_11;
input 	dffe121;
input 	dffe13;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	dffe101;
input 	dffe111;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~3 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \xordvalue~0_combout ;


NCO_Lab3_lpm_add_sub_22 u0(
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.dffe12(dffe12),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe13),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout(\Add0~3 ));
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(\Add0~3 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000000000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_22 (
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	a_0,
	xordvalue_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg_8 auto_generated(
	.dffe13(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.dffe121(dffe12),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg_8 (
	dffe13,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	a_0,
	xordvalue_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe13;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
output 	dffe111;
output 	dffe121;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;


dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm_9 (
	dffe12,
	a_0,
	xordvalue_2,
	dffe16,
	cor1x_10,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe1,
	dffe2,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
input 	a_0;
input 	xordvalue_2;
input 	dffe16;
input 	cor1x_10;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe1;
output 	dffe2;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[11]~q ;
wire \Add0~0_combout ;
wire \a[10]~q ;
wire \Add0~1_combout ;


NCO_Lab3_lpm_add_sub_23 u0(
	.dffe12(dffe12),
	.a_0(a_0),
	.xordvalue_2(xordvalue_2),
	.a_11(\a[11]~q ),
	.dffe11(dffe11),
	.a_10(\a[10]~q ),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

cyclonev_lcell_comb \Add0~0 (
	.dataa(!dffe16),
	.datab(!cor1x_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Add0~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(!dffe16),
	.datab(!cor1x_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h7777777777777777;
defparam \Add0~1 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_23 (
	dffe12,
	a_0,
	xordvalue_2,
	a_11,
	dffe11,
	a_10,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe1,
	dffe2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
input 	a_0;
input 	xordvalue_2;
input 	a_11;
output 	dffe11;
input 	a_10;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe1;
output 	dffe2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg_9 auto_generated(
	.dffe121(dffe12),
	.a_0(a_0),
	.xordvalue_2(xordvalue_2),
	.a_11(a_11),
	.dffe111(dffe11),
	.a_10(a_10),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe13(dffe1),
	.dffe21(dffe2),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg_9 (
	dffe121,
	a_0,
	xordvalue_2,
	a_11,
	dffe111,
	a_10,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe13,
	dffe21,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe121;
input 	a_0;
input 	xordvalue_2;
input 	a_11;
output 	dffe111;
input 	a_10;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe13;
output 	dffe21;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;


dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!xordvalue_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_sxor_1p_lpm_10 (
	dffe12,
	dffe11,
	dffe16,
	dffe10,
	pipeline_dffe_11,
	dffe121,
	dffe9,
	pipeline_dffe_10,
	dffe8,
	pipeline_dffe_9,
	dffe111,
	dffe7,
	pipeline_dffe_8,
	dffe101,
	dffe6,
	pipeline_dffe_7,
	dffe91,
	dffe5,
	pipeline_dffe_6,
	dffe81,
	dffe4,
	dffe1,
	pipeline_dffe_5,
	dffe71,
	dffe2,
	dffe3,
	pipeline_dffe_4,
	dffe61,
	pipeline_dffe_3,
	dffe51,
	pipeline_dffe_2,
	dffe41,
	dffe31,
	dffe13,
	dffe21,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
input 	dffe16;
output 	dffe10;
input 	pipeline_dffe_11;
input 	dffe121;
output 	dffe9;
input 	pipeline_dffe_10;
output 	dffe8;
input 	pipeline_dffe_9;
input 	dffe111;
output 	dffe7;
input 	pipeline_dffe_8;
input 	dffe101;
output 	dffe6;
input 	pipeline_dffe_7;
input 	dffe91;
output 	dffe5;
input 	pipeline_dffe_6;
input 	dffe81;
output 	dffe4;
output 	dffe1;
input 	pipeline_dffe_5;
input 	dffe71;
output 	dffe2;
output 	dffe3;
input 	pipeline_dffe_4;
input 	dffe61;
input 	pipeline_dffe_3;
input 	dffe51;
input 	pipeline_dffe_2;
input 	dffe41;
input 	dffe31;
input 	dffe13;
input 	dffe21;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[11]~q ;
wire \xordvalue[10]~q ;
wire \xordvalue~0_combout ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \xordvalue~1_combout ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \xordvalue~2_combout ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \xordvalue~3_combout ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \xordvalue~4_combout ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \xordvalue~5_combout ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \xordvalue~6_combout ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;


NCO_Lab3_lpm_add_sub_24 u0(
	.dffe12(dffe12),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.dffe4(dffe4),
	.dffe1(dffe1),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe13),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

cyclonev_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

cyclonev_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

cyclonev_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

cyclonev_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

cyclonev_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

cyclonev_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

cyclonev_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

cyclonev_lcell_comb \xordvalue~9 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_24 (
	dffe12,
	dffe11,
	a_11,
	xordvalue_10,
	dffe10,
	a_10,
	dffe9,
	a_9,
	dffe8,
	a_8,
	xordvalue_8,
	dffe7,
	a_7,
	xordvalue_7,
	dffe6,
	a_6,
	xordvalue_6,
	dffe5,
	a_5,
	xordvalue_5,
	dffe4,
	dffe1,
	a_4,
	xordvalue_4,
	dffe2,
	dffe3,
	a_3,
	xordvalue_3,
	a_0,
	xordvalue_0,
	a_2,
	xordvalue_2,
	a_1,
	xordvalue_1,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe12;
output 	dffe11;
input 	a_11;
input 	xordvalue_10;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
input 	a_8;
input 	xordvalue_8;
output 	dffe7;
input 	a_7;
input 	xordvalue_7;
output 	dffe6;
input 	a_6;
input 	xordvalue_6;
output 	dffe5;
input 	a_5;
input 	xordvalue_5;
output 	dffe4;
output 	dffe1;
input 	a_4;
input 	xordvalue_4;
output 	dffe2;
output 	dffe3;
input 	a_3;
input 	xordvalue_3;
input 	a_0;
input 	xordvalue_0;
input 	a_2;
input 	xordvalue_2;
input 	a_1;
input 	xordvalue_1;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_bkg_10 auto_generated(
	.dffe121(dffe12),
	.dffe111(dffe11),
	.a_11(a_11),
	.xordvalue_10(xordvalue_10),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.dffe71(dffe7),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.dffe61(dffe6),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.dffe51(dffe5),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.dffe41(dffe4),
	.dffe13(dffe1),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_bkg_10 (
	dffe121,
	dffe111,
	a_11,
	xordvalue_10,
	dffe101,
	a_10,
	dffe91,
	a_9,
	dffe81,
	a_8,
	xordvalue_8,
	dffe71,
	a_7,
	xordvalue_7,
	dffe61,
	a_6,
	xordvalue_6,
	dffe51,
	a_5,
	xordvalue_5,
	dffe41,
	dffe13,
	a_4,
	xordvalue_4,
	dffe21,
	dffe31,
	a_3,
	xordvalue_3,
	a_0,
	xordvalue_0,
	a_2,
	xordvalue_2,
	a_1,
	xordvalue_1,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe121;
output 	dffe111;
input 	a_11;
input 	xordvalue_10;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
input 	a_8;
input 	xordvalue_8;
output 	dffe71;
input 	a_7;
input 	xordvalue_7;
output 	dffe61;
input 	a_6;
input 	xordvalue_6;
output 	dffe51;
input 	a_5;
input 	xordvalue_5;
output 	dffe41;
output 	dffe13;
input 	a_4;
input 	xordvalue_4;
output 	dffe21;
output 	dffe31;
input 	a_3;
input 	xordvalue_3;
input 	a_0;
input 	xordvalue_0;
input 	a_2;
input 	xordvalue_2;
input 	a_1;
input 	xordvalue_1;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;


dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe13),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm (
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \xordvalue[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \xordvalue[11]~0_combout ;


NCO_Lab3_lpm_add_sub_25 u0(
	.dffe16(dffe16),
	.dffe15(dffe15),
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.dffe14(dffe14),
	.a_14(\a[14]~q ),
	.dffe13(dffe13),
	.a_13(\a[13]~q ),
	.dffe12(dffe12),
	.a_12(\a[12]~q ),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.dffe4(dffe4),
	.a_4(\a[4]~q ),
	.dffe3(dffe3),
	.a_3(\a[3]~q ),
	.dffe2(dffe2),
	.a_2(\a[2]~q ),
	.dffe1(dffe1),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue[11]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue[11]~0 (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue[11]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue[11]~0 .extended_lut = "off";
defparam \xordvalue[11]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \xordvalue[11]~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_25 (
	dffe16,
	dffe15,
	a_15,
	xordvalue_0,
	dffe14,
	a_14,
	dffe13,
	a_13,
	dffe12,
	a_12,
	dffe11,
	a_11,
	xordvalue_11,
	dffe10,
	a_10,
	dffe9,
	a_9,
	dffe8,
	a_8,
	dffe7,
	a_7,
	dffe6,
	a_6,
	dffe5,
	a_5,
	dffe4,
	a_4,
	dffe3,
	a_3,
	dffe2,
	a_2,
	dffe1,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
input 	a_15;
input 	xordvalue_0;
output 	dffe14;
input 	a_14;
output 	dffe13;
input 	a_13;
output 	dffe12;
input 	a_12;
output 	dffe11;
input 	a_11;
input 	xordvalue_11;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
input 	a_8;
output 	dffe7;
input 	a_7;
output 	dffe6;
input 	a_6;
output 	dffe5;
input 	a_5;
output 	dffe4;
input 	a_4;
output 	dffe3;
input 	a_3;
output 	dffe2;
input 	a_2;
output 	dffe1;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg auto_generated(
	.dffe161(dffe16),
	.dffe151(dffe15),
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.dffe141(dffe14),
	.a_14(a_14),
	.dffe131(dffe13),
	.a_13(a_13),
	.dffe121(dffe12),
	.a_12(a_12),
	.dffe111(dffe11),
	.a_11(a_11),
	.xordvalue_11(xordvalue_11),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.a_8(a_8),
	.dffe71(dffe7),
	.a_7(a_7),
	.dffe61(dffe6),
	.a_6(a_6),
	.dffe51(dffe5),
	.a_5(a_5),
	.dffe41(dffe4),
	.a_4(a_4),
	.dffe31(dffe3),
	.a_3(a_3),
	.dffe21(dffe2),
	.a_2(a_2),
	.dffe17(dffe1),
	.a_1(a_1),
	.a_0(a_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg (
	dffe161,
	dffe151,
	a_15,
	xordvalue_0,
	dffe141,
	a_14,
	dffe131,
	a_13,
	dffe121,
	a_12,
	dffe111,
	a_11,
	xordvalue_11,
	dffe101,
	a_10,
	dffe91,
	a_9,
	dffe81,
	a_8,
	dffe71,
	a_7,
	dffe61,
	a_6,
	dffe51,
	a_5,
	dffe41,
	a_4,
	dffe31,
	a_3,
	dffe21,
	a_2,
	dffe17,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
output 	dffe151;
input 	a_15;
input 	xordvalue_0;
output 	dffe141;
input 	a_14;
output 	dffe131;
input 	a_13;
output 	dffe121;
input 	a_12;
output 	dffe111;
input 	a_11;
input 	xordvalue_11;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
input 	a_8;
output 	dffe71;
input 	a_7;
output 	dffe61;
input 	a_6;
output 	dffe51;
input 	a_5;
output 	dffe41;
input 	a_4;
output 	dffe31;
input 	a_3;
output 	dffe21;
input 	a_2;
output 	dffe17;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm_1 (
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \xordvalue[10]~0_combout ;


NCO_Lab3_lpm_add_sub_26 u0(
	.dffe16(dffe16),
	.dffe15(dffe15),
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.dffe14(dffe14),
	.a_14(\a[14]~q ),
	.dffe13(dffe13),
	.a_13(\a[13]~q ),
	.dffe12(dffe12),
	.a_12(\a[12]~q ),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.dffe4(dffe4),
	.a_4(\a[4]~q ),
	.dffe3(dffe3),
	.a_3(\a[3]~q ),
	.dffe2(dffe2),
	.a_2(\a[2]~q ),
	.dffe1(dffe1),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue[10]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue[10]~0 (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue[10]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue[10]~0 .extended_lut = "off";
defparam \xordvalue[10]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \xordvalue[10]~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_26 (
	dffe16,
	dffe15,
	a_15,
	xordvalue_0,
	dffe14,
	a_14,
	dffe13,
	a_13,
	dffe12,
	a_12,
	dffe11,
	a_11,
	dffe10,
	a_10,
	xordvalue_10,
	dffe9,
	a_9,
	dffe8,
	a_8,
	dffe7,
	a_7,
	dffe6,
	a_6,
	dffe5,
	a_5,
	dffe4,
	a_4,
	dffe3,
	a_3,
	dffe2,
	a_2,
	dffe1,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
input 	a_15;
input 	xordvalue_0;
output 	dffe14;
input 	a_14;
output 	dffe13;
input 	a_13;
output 	dffe12;
input 	a_12;
output 	dffe11;
input 	a_11;
output 	dffe10;
input 	a_10;
input 	xordvalue_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
input 	a_8;
output 	dffe7;
input 	a_7;
output 	dffe6;
input 	a_6;
output 	dffe5;
input 	a_5;
output 	dffe4;
input 	a_4;
output 	dffe3;
input 	a_3;
output 	dffe2;
input 	a_2;
output 	dffe1;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg_1 auto_generated(
	.dffe161(dffe16),
	.dffe151(dffe15),
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.dffe141(dffe14),
	.a_14(a_14),
	.dffe131(dffe13),
	.a_13(a_13),
	.dffe121(dffe12),
	.a_12(a_12),
	.dffe111(dffe11),
	.a_11(a_11),
	.dffe101(dffe10),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.a_8(a_8),
	.dffe71(dffe7),
	.a_7(a_7),
	.dffe61(dffe6),
	.a_6(a_6),
	.dffe51(dffe5),
	.a_5(a_5),
	.dffe41(dffe4),
	.a_4(a_4),
	.dffe31(dffe3),
	.a_3(a_3),
	.dffe21(dffe2),
	.a_2(a_2),
	.dffe17(dffe1),
	.a_1(a_1),
	.a_0(a_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg_1 (
	dffe161,
	dffe151,
	a_15,
	xordvalue_0,
	dffe141,
	a_14,
	dffe131,
	a_13,
	dffe121,
	a_12,
	dffe111,
	a_11,
	dffe101,
	a_10,
	xordvalue_10,
	dffe91,
	a_9,
	dffe81,
	a_8,
	dffe71,
	a_7,
	dffe61,
	a_6,
	dffe51,
	a_5,
	dffe41,
	a_4,
	dffe31,
	a_3,
	dffe21,
	a_2,
	dffe17,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
output 	dffe151;
input 	a_15;
input 	xordvalue_0;
output 	dffe141;
input 	a_14;
output 	dffe131;
input 	a_13;
output 	dffe121;
input 	a_12;
output 	dffe111;
input 	a_11;
output 	dffe101;
input 	a_10;
input 	xordvalue_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
input 	a_8;
output 	dffe71;
input 	a_7;
output 	dffe61;
input 	a_6;
output 	dffe51;
input 	a_5;
output 	dffe41;
input 	a_4;
output 	dffe31;
input 	a_3;
output 	dffe21;
input 	a_2;
output 	dffe17;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm_2 (
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \a[15]~q ;
wire \xordvalue[10]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \xordvalue[0]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~0_combout ;


NCO_Lab3_lpm_add_sub_27 u0(
	.dffe16(dffe16),
	.dffe15(dffe15),
	.a_15(\a[15]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe14(dffe14),
	.a_14(\a[14]~q ),
	.dffe13(dffe13),
	.a_13(\a[13]~q ),
	.dffe12(dffe12),
	.a_12(\a[12]~q ),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.dffe4(dffe4),
	.a_4(\a[4]~q ),
	.dffe3(dffe3),
	.a_3(\a[3]~q ),
	.dffe2(dffe2),
	.a_2(\a[2]~q ),
	.dffe1(dffe1),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue[0]~0 (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue[0]~0 .extended_lut = "off";
defparam \xordvalue[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \xordvalue[0]~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_27 (
	dffe16,
	dffe15,
	a_15,
	xordvalue_10,
	dffe14,
	a_14,
	dffe13,
	a_13,
	dffe12,
	a_12,
	dffe11,
	a_11,
	dffe10,
	a_10,
	dffe9,
	a_9,
	xordvalue_0,
	dffe8,
	a_8,
	dffe7,
	a_7,
	dffe6,
	a_6,
	dffe5,
	a_5,
	dffe4,
	a_4,
	dffe3,
	a_3,
	dffe2,
	a_2,
	dffe1,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
input 	a_15;
input 	xordvalue_10;
output 	dffe14;
input 	a_14;
output 	dffe13;
input 	a_13;
output 	dffe12;
input 	a_12;
output 	dffe11;
input 	a_11;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
input 	xordvalue_0;
output 	dffe8;
input 	a_8;
output 	dffe7;
input 	a_7;
output 	dffe6;
input 	a_6;
output 	dffe5;
input 	a_5;
output 	dffe4;
input 	a_4;
output 	dffe3;
input 	a_3;
output 	dffe2;
input 	a_2;
output 	dffe1;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg_2 auto_generated(
	.dffe161(dffe16),
	.dffe151(dffe15),
	.a_15(a_15),
	.xordvalue_10(xordvalue_10),
	.dffe141(dffe14),
	.a_14(a_14),
	.dffe131(dffe13),
	.a_13(a_13),
	.dffe121(dffe12),
	.a_12(a_12),
	.dffe111(dffe11),
	.a_11(a_11),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.xordvalue_0(xordvalue_0),
	.dffe81(dffe8),
	.a_8(a_8),
	.dffe71(dffe7),
	.a_7(a_7),
	.dffe61(dffe6),
	.a_6(a_6),
	.dffe51(dffe5),
	.a_5(a_5),
	.dffe41(dffe4),
	.a_4(a_4),
	.dffe31(dffe3),
	.a_3(a_3),
	.dffe21(dffe2),
	.a_2(a_2),
	.dffe17(dffe1),
	.a_1(a_1),
	.a_0(a_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg_2 (
	dffe161,
	dffe151,
	a_15,
	xordvalue_10,
	dffe141,
	a_14,
	dffe131,
	a_13,
	dffe121,
	a_12,
	dffe111,
	a_11,
	dffe101,
	a_10,
	dffe91,
	a_9,
	xordvalue_0,
	dffe81,
	a_8,
	dffe71,
	a_7,
	dffe61,
	a_6,
	dffe51,
	a_5,
	dffe41,
	a_4,
	dffe31,
	a_3,
	dffe21,
	a_2,
	dffe17,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
output 	dffe151;
input 	a_15;
input 	xordvalue_10;
output 	dffe141;
input 	a_14;
output 	dffe131;
input 	a_13;
output 	dffe121;
input 	a_12;
output 	dffe111;
input 	a_11;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
input 	xordvalue_0;
output 	dffe81;
input 	a_8;
output 	dffe71;
input 	a_7;
output 	dffe61;
input 	a_6;
output 	dffe51;
input 	a_5;
output 	dffe41;
input 	a_4;
output 	dffe31;
input 	a_3;
output 	dffe21;
input 	a_2;
output 	dffe17;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm_3 (
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \a[15]~q ;
wire \xordvalue[10]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \xordvalue[0]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~0_combout ;


NCO_Lab3_lpm_add_sub_28 u0(
	.dffe16(dffe16),
	.dffe15(dffe15),
	.a_15(\a[15]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe14(dffe14),
	.a_14(\a[14]~q ),
	.dffe13(dffe13),
	.a_13(\a[13]~q ),
	.dffe12(dffe12),
	.a_12(\a[12]~q ),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.dffe4(dffe4),
	.a_4(\a[4]~q ),
	.dffe3(dffe3),
	.a_3(\a[3]~q ),
	.dffe2(dffe2),
	.a_2(\a[2]~q ),
	.dffe1(dffe1),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue[0]~0 (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue[0]~0 .extended_lut = "off";
defparam \xordvalue[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \xordvalue[0]~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_28 (
	dffe16,
	dffe15,
	a_15,
	xordvalue_10,
	dffe14,
	a_14,
	dffe13,
	a_13,
	dffe12,
	a_12,
	dffe11,
	a_11,
	dffe10,
	a_10,
	dffe9,
	a_9,
	dffe8,
	a_8,
	xordvalue_0,
	dffe7,
	a_7,
	dffe6,
	a_6,
	dffe5,
	a_5,
	dffe4,
	a_4,
	dffe3,
	a_3,
	dffe2,
	a_2,
	dffe1,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
input 	a_15;
input 	xordvalue_10;
output 	dffe14;
input 	a_14;
output 	dffe13;
input 	a_13;
output 	dffe12;
input 	a_12;
output 	dffe11;
input 	a_11;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
input 	a_8;
input 	xordvalue_0;
output 	dffe7;
input 	a_7;
output 	dffe6;
input 	a_6;
output 	dffe5;
input 	a_5;
output 	dffe4;
input 	a_4;
output 	dffe3;
input 	a_3;
output 	dffe2;
input 	a_2;
output 	dffe1;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg_3 auto_generated(
	.dffe161(dffe16),
	.dffe151(dffe15),
	.a_15(a_15),
	.xordvalue_10(xordvalue_10),
	.dffe141(dffe14),
	.a_14(a_14),
	.dffe131(dffe13),
	.a_13(a_13),
	.dffe121(dffe12),
	.a_12(a_12),
	.dffe111(dffe11),
	.a_11(a_11),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.a_8(a_8),
	.xordvalue_0(xordvalue_0),
	.dffe71(dffe7),
	.a_7(a_7),
	.dffe61(dffe6),
	.a_6(a_6),
	.dffe51(dffe5),
	.a_5(a_5),
	.dffe41(dffe4),
	.a_4(a_4),
	.dffe31(dffe3),
	.a_3(a_3),
	.dffe21(dffe2),
	.a_2(a_2),
	.dffe17(dffe1),
	.a_1(a_1),
	.a_0(a_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg_3 (
	dffe161,
	dffe151,
	a_15,
	xordvalue_10,
	dffe141,
	a_14,
	dffe131,
	a_13,
	dffe121,
	a_12,
	dffe111,
	a_11,
	dffe101,
	a_10,
	dffe91,
	a_9,
	dffe81,
	a_8,
	xordvalue_0,
	dffe71,
	a_7,
	dffe61,
	a_6,
	dffe51,
	a_5,
	dffe41,
	a_4,
	dffe31,
	a_3,
	dffe21,
	a_2,
	dffe17,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
output 	dffe151;
input 	a_15;
input 	xordvalue_10;
output 	dffe141;
input 	a_14;
output 	dffe131;
input 	a_13;
output 	dffe121;
input 	a_12;
output 	dffe111;
input 	a_11;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
input 	a_8;
input 	xordvalue_0;
output 	dffe71;
input 	a_7;
output 	dffe61;
input 	a_6;
output 	dffe51;
input 	a_5;
output 	dffe41;
input 	a_4;
output 	dffe31;
input 	a_3;
output 	dffe21;
input 	a_2;
output 	dffe17;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm_4 (
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \xordvalue[1]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \xordvalue[1]~0_combout ;


NCO_Lab3_lpm_add_sub_29 u0(
	.dffe16(dffe16),
	.dffe15(dffe15),
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.dffe14(dffe14),
	.a_14(\a[14]~q ),
	.dffe13(dffe13),
	.a_13(\a[13]~q ),
	.dffe12(dffe12),
	.a_12(\a[12]~q ),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.dffe4(dffe4),
	.a_4(\a[4]~q ),
	.dffe3(dffe3),
	.a_3(\a[3]~q ),
	.dffe2(dffe2),
	.a_2(\a[2]~q ),
	.dffe1(dffe1),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue[1]~0 (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue[1]~0 .extended_lut = "off";
defparam \xordvalue[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \xordvalue[1]~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_29 (
	dffe16,
	dffe15,
	a_15,
	xordvalue_0,
	dffe14,
	a_14,
	dffe13,
	a_13,
	dffe12,
	a_12,
	dffe11,
	a_11,
	dffe10,
	a_10,
	dffe9,
	a_9,
	dffe8,
	a_8,
	dffe7,
	a_7,
	xordvalue_1,
	dffe6,
	a_6,
	dffe5,
	a_5,
	dffe4,
	a_4,
	dffe3,
	a_3,
	dffe2,
	a_2,
	dffe1,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
input 	a_15;
input 	xordvalue_0;
output 	dffe14;
input 	a_14;
output 	dffe13;
input 	a_13;
output 	dffe12;
input 	a_12;
output 	dffe11;
input 	a_11;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
input 	a_8;
output 	dffe7;
input 	a_7;
input 	xordvalue_1;
output 	dffe6;
input 	a_6;
output 	dffe5;
input 	a_5;
output 	dffe4;
input 	a_4;
output 	dffe3;
input 	a_3;
output 	dffe2;
input 	a_2;
output 	dffe1;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg_4 auto_generated(
	.dffe161(dffe16),
	.dffe151(dffe15),
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.dffe141(dffe14),
	.a_14(a_14),
	.dffe131(dffe13),
	.a_13(a_13),
	.dffe121(dffe12),
	.a_12(a_12),
	.dffe111(dffe11),
	.a_11(a_11),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.a_8(a_8),
	.dffe71(dffe7),
	.a_7(a_7),
	.xordvalue_1(xordvalue_1),
	.dffe61(dffe6),
	.a_6(a_6),
	.dffe51(dffe5),
	.a_5(a_5),
	.dffe41(dffe4),
	.a_4(a_4),
	.dffe31(dffe3),
	.a_3(a_3),
	.dffe21(dffe2),
	.a_2(a_2),
	.dffe17(dffe1),
	.a_1(a_1),
	.a_0(a_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg_4 (
	dffe161,
	dffe151,
	a_15,
	xordvalue_0,
	dffe141,
	a_14,
	dffe131,
	a_13,
	dffe121,
	a_12,
	dffe111,
	a_11,
	dffe101,
	a_10,
	dffe91,
	a_9,
	dffe81,
	a_8,
	dffe71,
	a_7,
	xordvalue_1,
	dffe61,
	a_6,
	dffe51,
	a_5,
	dffe41,
	a_4,
	dffe31,
	a_3,
	dffe21,
	a_2,
	dffe17,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
output 	dffe151;
input 	a_15;
input 	xordvalue_0;
output 	dffe141;
input 	a_14;
output 	dffe131;
input 	a_13;
output 	dffe121;
input 	a_12;
output 	dffe111;
input 	a_11;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
input 	a_8;
output 	dffe71;
input 	a_7;
input 	xordvalue_1;
output 	dffe61;
input 	a_6;
output 	dffe51;
input 	a_5;
output 	dffe41;
input 	a_4;
output 	dffe31;
input 	a_3;
output 	dffe21;
input 	a_2;
output 	dffe17;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm_5 (
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \a[15]~q ;
wire \xordvalue[10]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \xordvalue[0]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~0_combout ;


NCO_Lab3_lpm_add_sub_30 u0(
	.dffe16(dffe16),
	.dffe15(dffe15),
	.a_15(\a[15]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe14(dffe14),
	.a_14(\a[14]~q ),
	.dffe13(dffe13),
	.a_13(\a[13]~q ),
	.dffe12(dffe12),
	.a_12(\a[12]~q ),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.dffe4(dffe4),
	.a_4(\a[4]~q ),
	.dffe3(dffe3),
	.a_3(\a[3]~q ),
	.dffe2(dffe2),
	.a_2(\a[2]~q ),
	.dffe1(dffe1),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue[0]~0 (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue[0]~0 .extended_lut = "off";
defparam \xordvalue[0]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \xordvalue[0]~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_30 (
	dffe16,
	dffe15,
	a_15,
	xordvalue_10,
	dffe14,
	a_14,
	dffe13,
	a_13,
	dffe12,
	a_12,
	dffe11,
	a_11,
	dffe10,
	a_10,
	dffe9,
	a_9,
	dffe8,
	a_8,
	dffe7,
	a_7,
	dffe6,
	a_6,
	xordvalue_0,
	dffe5,
	a_5,
	dffe4,
	a_4,
	dffe3,
	a_3,
	dffe2,
	a_2,
	dffe1,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
input 	a_15;
input 	xordvalue_10;
output 	dffe14;
input 	a_14;
output 	dffe13;
input 	a_13;
output 	dffe12;
input 	a_12;
output 	dffe11;
input 	a_11;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
input 	a_8;
output 	dffe7;
input 	a_7;
output 	dffe6;
input 	a_6;
input 	xordvalue_0;
output 	dffe5;
input 	a_5;
output 	dffe4;
input 	a_4;
output 	dffe3;
input 	a_3;
output 	dffe2;
input 	a_2;
output 	dffe1;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg_5 auto_generated(
	.dffe161(dffe16),
	.dffe151(dffe15),
	.a_15(a_15),
	.xordvalue_10(xordvalue_10),
	.dffe141(dffe14),
	.a_14(a_14),
	.dffe131(dffe13),
	.a_13(a_13),
	.dffe121(dffe12),
	.a_12(a_12),
	.dffe111(dffe11),
	.a_11(a_11),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.a_8(a_8),
	.dffe71(dffe7),
	.a_7(a_7),
	.dffe61(dffe6),
	.a_6(a_6),
	.xordvalue_0(xordvalue_0),
	.dffe51(dffe5),
	.a_5(a_5),
	.dffe41(dffe4),
	.a_4(a_4),
	.dffe31(dffe3),
	.a_3(a_3),
	.dffe21(dffe2),
	.a_2(a_2),
	.dffe17(dffe1),
	.a_1(a_1),
	.a_0(a_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg_5 (
	dffe161,
	dffe151,
	a_15,
	xordvalue_10,
	dffe141,
	a_14,
	dffe131,
	a_13,
	dffe121,
	a_12,
	dffe111,
	a_11,
	dffe101,
	a_10,
	dffe91,
	a_9,
	dffe81,
	a_8,
	dffe71,
	a_7,
	dffe61,
	a_6,
	xordvalue_0,
	dffe51,
	a_5,
	dffe41,
	a_4,
	dffe31,
	a_3,
	dffe21,
	a_2,
	dffe17,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
output 	dffe151;
input 	a_15;
input 	xordvalue_10;
output 	dffe141;
input 	a_14;
output 	dffe131;
input 	a_13;
output 	dffe121;
input 	a_12;
output 	dffe111;
input 	a_11;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
input 	a_8;
output 	dffe71;
input 	a_7;
output 	dffe61;
input 	a_6;
input 	xordvalue_0;
output 	dffe51;
input 	a_5;
output 	dffe41;
input 	a_4;
output 	dffe31;
input 	a_3;
output 	dffe21;
input 	a_2;
output 	dffe17;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm_6 (
	dffe16,
	corx_10,
	dffe15,
	dffe14,
	corz_14,
	dffe13,
	corz_13,
	dffe12,
	corz_12,
	dffe11,
	corz_11,
	dffe10,
	corz_10,
	dffe9,
	corz_9,
	dffe8,
	corz_8,
	dffe7,
	corz_7,
	dffe6,
	corz_6,
	dffe5,
	corz_5,
	dffe4,
	corz_4,
	dffe3,
	corz_3,
	dffe2,
	corz_2,
	dffe1,
	corz_1,
	corz_0,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
input 	corx_10;
output 	dffe15;
output 	dffe14;
input 	corz_14;
output 	dffe13;
input 	corz_13;
output 	dffe12;
input 	corz_12;
output 	dffe11;
input 	corz_11;
output 	dffe10;
input 	corz_10;
output 	dffe9;
input 	corz_9;
output 	dffe8;
input 	corz_8;
output 	dffe7;
input 	corz_7;
output 	dffe6;
input 	corz_6;
output 	dffe5;
input 	corz_5;
output 	dffe4;
input 	corz_4;
output 	dffe3;
input 	corz_3;
output 	dffe2;
input 	corz_2;
output 	dffe1;
input 	corz_1;
input 	corz_0;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;


NCO_Lab3_lpm_add_sub_33 u0(
	.dffe16(dffe16),
	.corx_10(corx_10),
	.dffe15(dffe15),
	.a_14(\a[14]~q ),
	.dffe14(dffe14),
	.a_13(\a[13]~q ),
	.dffe13(dffe13),
	.a_12(\a[12]~q ),
	.dffe12(dffe12),
	.a_11(\a[11]~q ),
	.dffe11(dffe11),
	.a_10(\a[10]~q ),
	.dffe10(dffe10),
	.a_9(\a[9]~q ),
	.dffe9(dffe9),
	.a_8(\a[8]~q ),
	.dffe8(dffe8),
	.a_7(\a[7]~q ),
	.dffe7(dffe7),
	.a_6(\a[6]~q ),
	.dffe6(dffe6),
	.a_5(\a[5]~q ),
	.dffe5(dffe5),
	.a_4(\a[4]~q ),
	.dffe4(dffe4),
	.a_3(\a[3]~q ),
	.dffe3(dffe3),
	.a_2(\a[2]~q ),
	.dffe2(dffe2),
	.a_1(\a[1]~q ),
	.dffe1(dffe1),
	.a_0(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[14] (
	.clk(clk),
	.d(corz_14),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(corz_13),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(corz_12),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(corz_11),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(corz_10),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(corz_9),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(corz_8),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(corz_7),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(corz_6),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(corz_5),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(corz_4),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(corz_3),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(corz_2),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(corz_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(corz_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm_7 (
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \xordvalue[3]~0_combout ;


NCO_Lab3_lpm_add_sub_31 u0(
	.dffe16(dffe16),
	.dffe15(dffe15),
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.dffe14(dffe14),
	.a_14(\a[14]~q ),
	.dffe13(dffe13),
	.a_13(\a[13]~q ),
	.dffe12(dffe12),
	.a_12(\a[12]~q ),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.dffe4(dffe4),
	.a_4(\a[4]~q ),
	.dffe3(dffe3),
	.a_3(\a[3]~q ),
	.dffe2(dffe2),
	.a_2(\a[2]~q ),
	.dffe1(dffe1),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue[3]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue[3]~0 (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue[3]~0 .extended_lut = "off";
defparam \xordvalue[3]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \xordvalue[3]~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_31 (
	dffe16,
	dffe15,
	a_15,
	xordvalue_0,
	dffe14,
	a_14,
	dffe13,
	a_13,
	dffe12,
	a_12,
	dffe11,
	a_11,
	dffe10,
	a_10,
	dffe9,
	a_9,
	dffe8,
	a_8,
	dffe7,
	a_7,
	dffe6,
	a_6,
	dffe5,
	a_5,
	xordvalue_3,
	dffe4,
	a_4,
	dffe3,
	a_3,
	dffe2,
	a_2,
	dffe1,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
input 	a_15;
input 	xordvalue_0;
output 	dffe14;
input 	a_14;
output 	dffe13;
input 	a_13;
output 	dffe12;
input 	a_12;
output 	dffe11;
input 	a_11;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
input 	a_8;
output 	dffe7;
input 	a_7;
output 	dffe6;
input 	a_6;
output 	dffe5;
input 	a_5;
input 	xordvalue_3;
output 	dffe4;
input 	a_4;
output 	dffe3;
input 	a_3;
output 	dffe2;
input 	a_2;
output 	dffe1;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg_6 auto_generated(
	.dffe161(dffe16),
	.dffe151(dffe15),
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.dffe141(dffe14),
	.a_14(a_14),
	.dffe131(dffe13),
	.a_13(a_13),
	.dffe121(dffe12),
	.a_12(a_12),
	.dffe111(dffe11),
	.a_11(a_11),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.a_8(a_8),
	.dffe71(dffe7),
	.a_7(a_7),
	.dffe61(dffe6),
	.a_6(a_6),
	.dffe51(dffe5),
	.a_5(a_5),
	.xordvalue_3(xordvalue_3),
	.dffe41(dffe4),
	.a_4(a_4),
	.dffe31(dffe3),
	.a_3(a_3),
	.dffe21(dffe2),
	.a_2(a_2),
	.dffe17(dffe1),
	.a_1(a_1),
	.a_0(a_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg_6 (
	dffe161,
	dffe151,
	a_15,
	xordvalue_0,
	dffe141,
	a_14,
	dffe131,
	a_13,
	dffe121,
	a_12,
	dffe111,
	a_11,
	dffe101,
	a_10,
	dffe91,
	a_9,
	dffe81,
	a_8,
	dffe71,
	a_7,
	dffe61,
	a_6,
	dffe51,
	a_5,
	xordvalue_3,
	dffe41,
	a_4,
	dffe31,
	a_3,
	dffe21,
	a_2,
	dffe17,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
output 	dffe151;
input 	a_15;
input 	xordvalue_0;
output 	dffe141;
input 	a_14;
output 	dffe131;
input 	a_13;
output 	dffe121;
input 	a_12;
output 	dffe111;
input 	a_11;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
input 	a_8;
output 	dffe71;
input 	a_7;
output 	dffe61;
input 	a_6;
output 	dffe51;
input 	a_5;
input 	xordvalue_3;
output 	dffe41;
input 	a_4;
output 	dffe31;
input 	a_3;
output 	dffe21;
input 	a_2;
output 	dffe17;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm_8 (
	dffe16,
	dffe161,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
input 	dffe161;
input 	dffe15;
input 	dffe14;
input 	dffe13;
input 	dffe12;
input 	dffe11;
input 	dffe10;
input 	dffe9;
input 	dffe8;
input 	dffe7;
input 	dffe6;
input 	dffe5;
input 	dffe4;
input 	dffe3;
input 	dffe2;
input 	dffe1;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \xordvalue[2]~0_combout ;


NCO_Lab3_lpm_add_sub_32 u0(
	.dffe16(dffe16),
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe1),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue[2]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue[2]~0 (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue[2]~0 .extended_lut = "off";
defparam \xordvalue[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \xordvalue[2]~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_32 (
	dffe16,
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	xordvalue_2,
	a_3,
	a_2,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	xordvalue_2;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg_7 auto_generated(
	.dffe161(dffe16),
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg_7 (
	dffe161,
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	xordvalue_2,
	a_3,
	a_2,
	a_1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	xordvalue_2;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_33 (
	dffe16,
	corx_10,
	dffe15,
	a_14,
	dffe14,
	a_13,
	dffe13,
	a_12,
	dffe12,
	a_11,
	dffe11,
	a_10,
	dffe10,
	a_9,
	dffe9,
	a_8,
	dffe8,
	a_7,
	dffe7,
	a_6,
	dffe6,
	a_5,
	dffe5,
	a_4,
	dffe4,
	a_3,
	dffe3,
	a_2,
	dffe2,
	a_1,
	dffe1,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
input 	corx_10;
output 	dffe15;
input 	a_14;
output 	dffe14;
input 	a_13;
output 	dffe13;
input 	a_12;
output 	dffe12;
input 	a_11;
output 	dffe11;
input 	a_10;
output 	dffe10;
input 	a_9;
output 	dffe9;
input 	a_8;
output 	dffe8;
input 	a_7;
output 	dffe7;
input 	a_6;
output 	dffe6;
input 	a_5;
output 	dffe5;
input 	a_4;
output 	dffe4;
input 	a_3;
output 	dffe3;
input 	a_2;
output 	dffe2;
input 	a_1;
output 	dffe1;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg_8 auto_generated(
	.dffe161(dffe16),
	.corx_10(corx_10),
	.dffe151(dffe15),
	.a_14(a_14),
	.dffe141(dffe14),
	.a_13(a_13),
	.dffe131(dffe13),
	.a_12(a_12),
	.dffe121(dffe12),
	.a_11(a_11),
	.dffe111(dffe11),
	.a_10(a_10),
	.dffe101(dffe10),
	.a_9(a_9),
	.dffe91(dffe9),
	.a_8(a_8),
	.dffe81(dffe8),
	.a_7(a_7),
	.dffe71(dffe7),
	.a_6(a_6),
	.dffe61(dffe6),
	.a_5(a_5),
	.dffe51(dffe5),
	.a_4(a_4),
	.dffe41(dffe4),
	.a_3(a_3),
	.dffe31(dffe3),
	.a_2(a_2),
	.dffe21(dffe2),
	.a_1(a_1),
	.dffe17(dffe1),
	.a_0(a_0),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg_8 (
	dffe161,
	corx_10,
	dffe151,
	a_14,
	dffe141,
	a_13,
	dffe131,
	a_12,
	dffe121,
	a_11,
	dffe111,
	a_10,
	dffe101,
	a_9,
	dffe91,
	a_8,
	dffe81,
	a_7,
	dffe71,
	a_6,
	dffe61,
	a_5,
	dffe51,
	a_4,
	dffe41,
	a_3,
	dffe31,
	a_2,
	dffe21,
	a_1,
	dffe17,
	a_0,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
input 	corx_10;
output 	dffe151;
input 	a_14;
output 	dffe141;
input 	a_13;
output 	dffe131;
input 	a_12;
output 	dffe121;
input 	a_11;
output 	dffe111;
input 	a_10;
output 	dffe101;
input 	a_9;
output 	dffe91;
input 	a_8;
output 	dffe81;
input 	a_7;
output 	dffe71;
input 	a_6;
output 	dffe61;
input 	a_5;
output 	dffe51;
input 	a_4;
output 	dffe41;
input 	a_3;
output 	dffe31;
input 	a_2;
output 	dffe21;
input 	a_1;
output 	dffe17;
input 	a_0;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!corx_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm_9 (
	dffe16,
	a_0,
	dffe15,
	dffe161,
	dffe14,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
input 	a_0;
output 	dffe15;
input 	dffe161;
output 	dffe14;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \a[15]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \xordvalue[10]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \xordvalue[10]~0_combout ;


NCO_Lab3_lpm_add_sub_34 u0(
	.dffe16(dffe16),
	.a_0(a_0),
	.dffe15(dffe15),
	.a_15(\a[15]~q ),
	.dffe14(dffe14),
	.a_14(\a[14]~q ),
	.dffe13(dffe13),
	.a_13(\a[13]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.dffe12(dffe12),
	.a_12(\a[12]~q ),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.dffe4(dffe4),
	.a_4(\a[4]~q ),
	.dffe3(dffe3),
	.a_3(\a[3]~q ),
	.dffe2(dffe2),
	.a_2(\a[2]~q ),
	.dffe1(dffe1),
	.a_1(\a[1]~q ),
	.a_01(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue[10]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue[10]~0 (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue[10]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue[10]~0 .extended_lut = "off";
defparam \xordvalue[10]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \xordvalue[10]~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_34 (
	dffe16,
	a_0,
	dffe15,
	a_15,
	dffe14,
	a_14,
	dffe13,
	a_13,
	xordvalue_10,
	dffe12,
	a_12,
	dffe11,
	a_11,
	dffe10,
	a_10,
	dffe9,
	a_9,
	dffe8,
	a_8,
	dffe7,
	a_7,
	dffe6,
	a_6,
	dffe5,
	a_5,
	dffe4,
	a_4,
	dffe3,
	a_3,
	dffe2,
	a_2,
	dffe1,
	a_1,
	a_01,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
input 	a_0;
output 	dffe15;
input 	a_15;
output 	dffe14;
input 	a_14;
output 	dffe13;
input 	a_13;
input 	xordvalue_10;
output 	dffe12;
input 	a_12;
output 	dffe11;
input 	a_11;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
input 	a_8;
output 	dffe7;
input 	a_7;
output 	dffe6;
input 	a_6;
output 	dffe5;
input 	a_5;
output 	dffe4;
input 	a_4;
output 	dffe3;
input 	a_3;
output 	dffe2;
input 	a_2;
output 	dffe1;
input 	a_1;
input 	a_01;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg_9 auto_generated(
	.dffe161(dffe16),
	.a_0(a_0),
	.dffe151(dffe15),
	.a_15(a_15),
	.dffe141(dffe14),
	.a_14(a_14),
	.dffe131(dffe13),
	.a_13(a_13),
	.xordvalue_10(xordvalue_10),
	.dffe121(dffe12),
	.a_12(a_12),
	.dffe111(dffe11),
	.a_11(a_11),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.a_8(a_8),
	.dffe71(dffe7),
	.a_7(a_7),
	.dffe61(dffe6),
	.a_6(a_6),
	.dffe51(dffe5),
	.a_5(a_5),
	.dffe41(dffe4),
	.a_4(a_4),
	.dffe31(dffe3),
	.a_3(a_3),
	.dffe21(dffe2),
	.a_2(a_2),
	.dffe17(dffe1),
	.a_1(a_1),
	.a_01(a_01),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg_9 (
	dffe161,
	a_0,
	dffe151,
	a_15,
	dffe141,
	a_14,
	dffe131,
	a_13,
	xordvalue_10,
	dffe121,
	a_12,
	dffe111,
	a_11,
	dffe101,
	a_10,
	dffe91,
	a_9,
	dffe81,
	a_8,
	dffe71,
	a_7,
	dffe61,
	a_6,
	dffe51,
	a_5,
	dffe41,
	a_4,
	dffe31,
	a_3,
	dffe21,
	a_2,
	dffe17,
	a_1,
	a_01,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
input 	a_0;
output 	dffe151;
input 	a_15;
output 	dffe141;
input 	a_14;
output 	dffe131;
input 	a_13;
input 	xordvalue_10;
output 	dffe121;
input 	a_12;
output 	dffe111;
input 	a_11;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
input 	a_8;
output 	dffe71;
input 	a_7;
output 	dffe61;
input 	a_6;
output 	dffe51;
input 	a_5;
output 	dffe41;
input 	a_4;
output 	dffe31;
input 	a_3;
output 	dffe21;
input 	a_2;
output 	dffe17;
input 	a_1;
input 	a_01;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_01),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_cordic_zxor_1p_lpm_10 (
	dffe16,
	dffe15,
	a_0,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
input 	a_0;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \a[15]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \xordvalue[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \xordvalue[12]~0_combout ;


NCO_Lab3_lpm_add_sub_35 u0(
	.dffe16(dffe16),
	.dffe15(dffe15),
	.a_15(\a[15]~q ),
	.a_0(a_0),
	.dffe14(dffe14),
	.a_14(\a[14]~q ),
	.dffe13(dffe13),
	.a_13(\a[13]~q ),
	.dffe12(dffe12),
	.a_12(\a[12]~q ),
	.xordvalue_12(\xordvalue[12]~q ),
	.dffe11(dffe11),
	.a_11(\a[11]~q ),
	.dffe10(dffe10),
	.a_10(\a[10]~q ),
	.dffe9(dffe9),
	.a_9(\a[9]~q ),
	.dffe8(dffe8),
	.a_8(\a[8]~q ),
	.dffe7(dffe7),
	.a_7(\a[7]~q ),
	.dffe6(dffe6),
	.a_6(\a[6]~q ),
	.dffe5(dffe5),
	.a_5(\a[5]~q ),
	.dffe4(dffe4),
	.a_4(\a[4]~q ),
	.dffe3(dffe3),
	.a_3(\a[3]~q ),
	.dffe2(dffe2),
	.a_2(\a[2]~q ),
	.dffe1(dffe1),
	.a_1(\a[1]~q ),
	.a_01(\a[0]~q ),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \xordvalue[12] (
	.clk(clk),
	.d(\xordvalue[12]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\xordvalue[12]~q ),
	.prn(vcc));
defparam \xordvalue[12] .is_wysiwyg = "true";
defparam \xordvalue[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

cyclonev_lcell_comb \xordvalue[12]~0 (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue[12]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue[12]~0 .extended_lut = "off";
defparam \xordvalue[12]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \xordvalue[12]~0 .shared_arith = "off";

endmodule

module NCO_Lab3_lpm_add_sub_35 (
	dffe16,
	dffe15,
	a_15,
	a_0,
	dffe14,
	a_14,
	dffe13,
	a_13,
	dffe12,
	a_12,
	xordvalue_12,
	dffe11,
	a_11,
	dffe10,
	a_10,
	dffe9,
	a_9,
	dffe8,
	a_8,
	dffe7,
	a_7,
	dffe6,
	a_6,
	dffe5,
	a_5,
	dffe4,
	a_4,
	dffe3,
	a_3,
	dffe2,
	a_2,
	dffe1,
	a_1,
	a_01,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe16;
output 	dffe15;
input 	a_15;
input 	a_0;
output 	dffe14;
input 	a_14;
output 	dffe13;
input 	a_13;
output 	dffe12;
input 	a_12;
input 	xordvalue_12;
output 	dffe11;
input 	a_11;
output 	dffe10;
input 	a_10;
output 	dffe9;
input 	a_9;
output 	dffe8;
input 	a_8;
output 	dffe7;
input 	a_7;
output 	dffe6;
input 	a_6;
output 	dffe5;
input 	a_5;
output 	dffe4;
input 	a_4;
output 	dffe3;
input 	a_3;
output 	dffe2;
input 	a_2;
output 	dffe1;
input 	a_1;
input 	a_01;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



NCO_Lab3_add_sub_fkg_10 auto_generated(
	.dffe161(dffe16),
	.dffe151(dffe15),
	.a_15(a_15),
	.a_0(a_0),
	.dffe141(dffe14),
	.a_14(a_14),
	.dffe131(dffe13),
	.a_13(a_13),
	.dffe121(dffe12),
	.a_12(a_12),
	.xordvalue_12(xordvalue_12),
	.dffe111(dffe11),
	.a_11(a_11),
	.dffe101(dffe10),
	.a_10(a_10),
	.dffe91(dffe9),
	.a_9(a_9),
	.dffe81(dffe8),
	.a_8(a_8),
	.dffe71(dffe7),
	.a_7(a_7),
	.dffe61(dffe6),
	.a_6(a_6),
	.dffe51(dffe5),
	.a_5(a_5),
	.dffe41(dffe4),
	.a_4(a_4),
	.dffe31(dffe3),
	.a_3(a_3),
	.dffe21(dffe2),
	.a_2(a_2),
	.dffe17(dffe1),
	.a_1(a_1),
	.a_01(a_01),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module NCO_Lab3_add_sub_fkg_10 (
	dffe161,
	dffe151,
	a_15,
	a_0,
	dffe141,
	a_14,
	dffe131,
	a_13,
	dffe121,
	a_12,
	xordvalue_12,
	dffe111,
	a_11,
	dffe101,
	a_10,
	dffe91,
	a_9,
	dffe81,
	a_8,
	dffe71,
	a_7,
	dffe61,
	a_6,
	dffe51,
	a_5,
	dffe41,
	a_4,
	dffe31,
	a_3,
	dffe21,
	a_2,
	dffe17,
	a_1,
	a_01,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	dffe161;
output 	dffe151;
input 	a_15;
input 	a_0;
output 	dffe141;
input 	a_14;
output 	dffe131;
input 	a_13;
output 	dffe121;
input 	a_12;
input 	xordvalue_12;
output 	dffe111;
input 	a_11;
output 	dffe101;
input 	a_10;
output 	dffe91;
input 	a_9;
output 	dffe81;
input 	a_8;
output 	dffe71;
input 	a_7;
output 	dffe61;
input 	a_6;
output 	dffe51;
input 	a_5;
output 	dffe41;
input 	a_4;
output 	dffe31;
input 	a_3;
output 	dffe21;
input 	a_2;
output 	dffe17;
input 	a_1;
input 	a_01;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

cyclonev_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_01),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

cyclonev_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module NCO_Lab3_sop_reg (
	sin_o_0,
	sin_o_1,
	sin_o_2,
	sin_o_3,
	sin_o_4,
	sin_o_5,
	sin_o_6,
	sin_o_7,
	sin_o_8,
	sin_o_9,
	sin_o_10,
	sin_o_11,
	sin_o_01,
	sin_o_12,
	sin_o_21,
	sin_o_31,
	sin_o_41,
	sin_o_51,
	sin_o_61,
	sin_o_71,
	sin_o_81,
	sin_o_91,
	sin_o_101,
	sin_o_111,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	sin_o_0;
output 	sin_o_1;
output 	sin_o_2;
output 	sin_o_3;
output 	sin_o_4;
output 	sin_o_5;
output 	sin_o_6;
output 	sin_o_7;
output 	sin_o_8;
output 	sin_o_9;
output 	sin_o_10;
output 	sin_o_11;
input 	sin_o_01;
input 	sin_o_12;
input 	sin_o_21;
input 	sin_o_31;
input 	sin_o_41;
input 	sin_o_51;
input 	sin_o_61;
input 	sin_o_71;
input 	sin_o_81;
input 	sin_o_91;
input 	sin_o_101;
input 	sin_o_111;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \sin_o[0] (
	.clk(clk),
	.d(sin_o_01),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_0),
	.prn(vcc));
defparam \sin_o[0] .is_wysiwyg = "true";
defparam \sin_o[0] .power_up = "low";

dffeas \sin_o[1] (
	.clk(clk),
	.d(sin_o_12),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_1),
	.prn(vcc));
defparam \sin_o[1] .is_wysiwyg = "true";
defparam \sin_o[1] .power_up = "low";

dffeas \sin_o[2] (
	.clk(clk),
	.d(sin_o_21),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_2),
	.prn(vcc));
defparam \sin_o[2] .is_wysiwyg = "true";
defparam \sin_o[2] .power_up = "low";

dffeas \sin_o[3] (
	.clk(clk),
	.d(sin_o_31),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_3),
	.prn(vcc));
defparam \sin_o[3] .is_wysiwyg = "true";
defparam \sin_o[3] .power_up = "low";

dffeas \sin_o[4] (
	.clk(clk),
	.d(sin_o_41),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_4),
	.prn(vcc));
defparam \sin_o[4] .is_wysiwyg = "true";
defparam \sin_o[4] .power_up = "low";

dffeas \sin_o[5] (
	.clk(clk),
	.d(sin_o_51),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_5),
	.prn(vcc));
defparam \sin_o[5] .is_wysiwyg = "true";
defparam \sin_o[5] .power_up = "low";

dffeas \sin_o[6] (
	.clk(clk),
	.d(sin_o_61),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_6),
	.prn(vcc));
defparam \sin_o[6] .is_wysiwyg = "true";
defparam \sin_o[6] .power_up = "low";

dffeas \sin_o[7] (
	.clk(clk),
	.d(sin_o_71),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_7),
	.prn(vcc));
defparam \sin_o[7] .is_wysiwyg = "true";
defparam \sin_o[7] .power_up = "low";

dffeas \sin_o[8] (
	.clk(clk),
	.d(sin_o_81),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_8),
	.prn(vcc));
defparam \sin_o[8] .is_wysiwyg = "true";
defparam \sin_o[8] .power_up = "low";

dffeas \sin_o[9] (
	.clk(clk),
	.d(sin_o_91),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_9),
	.prn(vcc));
defparam \sin_o[9] .is_wysiwyg = "true";
defparam \sin_o[9] .power_up = "low";

dffeas \sin_o[10] (
	.clk(clk),
	.d(sin_o_101),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_10),
	.prn(vcc));
defparam \sin_o[10] .is_wysiwyg = "true";
defparam \sin_o[10] .power_up = "low";

dffeas \sin_o[11] (
	.clk(clk),
	.d(sin_o_111),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(sin_o_11),
	.prn(vcc));
defparam \sin_o[11] .is_wysiwyg = "true";
defparam \sin_o[11] .power_up = "low";

endmodule
